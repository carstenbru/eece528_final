// system.v

// Generated using ACDS version 15.0 145

`timescale 1 ps / 1 ps
module system (
		input  wire        alt_vip_itc_0_clocked_video_vid_clk,       // alt_vip_itc_0_clocked_video.vid_clk
		output wire [23:0] alt_vip_itc_0_clocked_video_vid_data,      //                            .vid_data
		output wire        alt_vip_itc_0_clocked_video_underflow,     //                            .underflow
		output wire        alt_vip_itc_0_clocked_video_vid_datavalid, //                            .vid_datavalid
		output wire        alt_vip_itc_0_clocked_video_vid_v_sync,    //                            .vid_v_sync
		output wire        alt_vip_itc_0_clocked_video_vid_h_sync,    //                            .vid_h_sync
		output wire        alt_vip_itc_0_clocked_video_vid_f,         //                            .vid_f
		output wire        alt_vip_itc_0_clocked_video_vid_h,         //                            .vid_h
		output wire        alt_vip_itc_0_clocked_video_vid_v,         //                            .vid_v
		input  wire [7:0]  analog1_x_export,                          //                   analog1_x.export
		input  wire [7:0]  analog1_y_export,                          //                   analog1_y.export
		input  wire [7:0]  analog2_x_export,                          //                   analog2_x.export
		input  wire [7:0]  analog2_y_export,                          //                   analog2_y.export
		input  wire        boton_a_export,                            //                     boton_a.export
		input  wire        boton_b_export,                            //                     boton_b.export
		input  wire        boton_down_export,                         //                  boton_down.export
		input  wire        boton_l_export,                            //                     boton_l.export
		input  wire        boton_left_export,                         //                  boton_left.export
		input  wire        boton_r_export,                            //                     boton_r.export
		input  wire        boton_right_export,                        //                 boton_right.export
		input  wire        boton_up_export,                           //                    boton_up.export
		input  wire        boton_x_export,                            //                     boton_x.export
		input  wire        boton_y_export,                            //                     boton_y.export
		input  wire        clk_clk,                                   //                         clk.clk
		output wire        epcs_dclk,                                 //                        epcs.dclk
		output wire        epcs_sce,                                  //                            .sce
		output wire        epcs_sdo,                                  //                            .sdo
		input  wire        epcs_data0,                                //                            .data0
		output wire [7:0]  pio_led_green_export,                      //               pio_led_green.export
		input  wire [3:0]  pio_sw_export,                             //                      pio_sw.export
		input  wire        reset_reset_n,                             //                       reset.reset_n
		output wire [12:0] sdram_addr,                                //                       sdram.addr
		output wire [1:0]  sdram_ba,                                  //                            .ba
		output wire        sdram_cas_n,                               //                            .cas_n
		output wire        sdram_cke,                                 //                            .cke
		output wire        sdram_cs_n,                                //                            .cs_n
		inout  wire [15:0] sdram_dq,                                  //                            .dq
		output wire [1:0]  sdram_dqm,                                 //                            .dqm
		output wire        sdram_ras_n,                               //                            .ras_n
		output wire        sdram_we_n,                                //                            .we_n
		input  wire        touch_panel_busy_export,                   //            touch_panel_busy.export
		input  wire        touch_panel_penirq_n_export,               //        touch_panel_penirq_n.export
		input  wire        touch_panel_spi_MISO,                      //             touch_panel_spi.MISO
		output wire        touch_panel_spi_MOSI,                      //                            .MOSI
		output wire        touch_panel_spi_SCLK,                      //                            .SCLK
		output wire        touch_panel_spi_SS_n                       //                            .SS_n
	);

	wire         alt_vip_vfr_0_avalon_streaming_source_valid;                   // alt_vip_vfr_0:dout_valid -> alt_vip_itc_0:is_valid
	wire  [23:0] alt_vip_vfr_0_avalon_streaming_source_data;                    // alt_vip_vfr_0:dout_data -> alt_vip_itc_0:is_data
	wire         alt_vip_vfr_0_avalon_streaming_source_ready;                   // alt_vip_itc_0:is_ready -> alt_vip_vfr_0:dout_ready
	wire         alt_vip_vfr_0_avalon_streaming_source_startofpacket;           // alt_vip_vfr_0:dout_startofpacket -> alt_vip_itc_0:is_sop
	wire         alt_vip_vfr_0_avalon_streaming_source_endofpacket;             // alt_vip_vfr_0:dout_endofpacket -> alt_vip_itc_0:is_eop
	wire  [31:0] alt_vip_vfr_0_avalon_master_readdata;                          // mm_interconnect_0:alt_vip_vfr_0_avalon_master_readdata -> alt_vip_vfr_0:master_readdata
	wire         alt_vip_vfr_0_avalon_master_waitrequest;                       // mm_interconnect_0:alt_vip_vfr_0_avalon_master_waitrequest -> alt_vip_vfr_0:master_waitrequest
	wire  [31:0] alt_vip_vfr_0_avalon_master_address;                           // alt_vip_vfr_0:master_address -> mm_interconnect_0:alt_vip_vfr_0_avalon_master_address
	wire         alt_vip_vfr_0_avalon_master_read;                              // alt_vip_vfr_0:master_read -> mm_interconnect_0:alt_vip_vfr_0_avalon_master_read
	wire         alt_vip_vfr_0_avalon_master_readdatavalid;                     // mm_interconnect_0:alt_vip_vfr_0_avalon_master_readdatavalid -> alt_vip_vfr_0:master_readdatavalid
	wire   [5:0] alt_vip_vfr_0_avalon_master_burstcount;                        // alt_vip_vfr_0:master_burstcount -> mm_interconnect_0:alt_vip_vfr_0_avalon_master_burstcount
	wire  [31:0] cpu_data_master_readdata;                                      // mm_interconnect_0:cpu_data_master_readdata -> cpu:d_readdata
	wire         cpu_data_master_waitrequest;                                   // mm_interconnect_0:cpu_data_master_waitrequest -> cpu:d_waitrequest
	wire         cpu_data_master_debugaccess;                                   // cpu:jtag_debug_module_debugaccess_to_roms -> mm_interconnect_0:cpu_data_master_debugaccess
	wire  [25:0] cpu_data_master_address;                                       // cpu:d_address -> mm_interconnect_0:cpu_data_master_address
	wire   [3:0] cpu_data_master_byteenable;                                    // cpu:d_byteenable -> mm_interconnect_0:cpu_data_master_byteenable
	wire         cpu_data_master_read;                                          // cpu:d_read -> mm_interconnect_0:cpu_data_master_read
	wire         cpu_data_master_write;                                         // cpu:d_write -> mm_interconnect_0:cpu_data_master_write
	wire  [31:0] cpu_data_master_writedata;                                     // cpu:d_writedata -> mm_interconnect_0:cpu_data_master_writedata
	wire  [31:0] cpu_instruction_master_readdata;                               // mm_interconnect_0:cpu_instruction_master_readdata -> cpu:i_readdata
	wire         cpu_instruction_master_waitrequest;                            // mm_interconnect_0:cpu_instruction_master_waitrequest -> cpu:i_waitrequest
	wire  [25:0] cpu_instruction_master_address;                                // cpu:i_address -> mm_interconnect_0:cpu_instruction_master_address
	wire         cpu_instruction_master_read;                                   // cpu:i_read -> mm_interconnect_0:cpu_instruction_master_read
	wire         cpu_instruction_master_readdatavalid;                          // mm_interconnect_0:cpu_instruction_master_readdatavalid -> cpu:i_readdatavalid
	wire         mm_interconnect_0_sdram_s1_chipselect;                         // mm_interconnect_0:sdram_s1_chipselect -> sdram:az_cs
	wire  [15:0] mm_interconnect_0_sdram_s1_readdata;                           // sdram:za_data -> mm_interconnect_0:sdram_s1_readdata
	wire         mm_interconnect_0_sdram_s1_waitrequest;                        // sdram:za_waitrequest -> mm_interconnect_0:sdram_s1_waitrequest
	wire  [23:0] mm_interconnect_0_sdram_s1_address;                            // mm_interconnect_0:sdram_s1_address -> sdram:az_addr
	wire         mm_interconnect_0_sdram_s1_read;                               // mm_interconnect_0:sdram_s1_read -> sdram:az_rd_n
	wire   [1:0] mm_interconnect_0_sdram_s1_byteenable;                         // mm_interconnect_0:sdram_s1_byteenable -> sdram:az_be_n
	wire         mm_interconnect_0_sdram_s1_readdatavalid;                      // sdram:za_valid -> mm_interconnect_0:sdram_s1_readdatavalid
	wire         mm_interconnect_0_sdram_s1_write;                              // mm_interconnect_0:sdram_s1_write -> sdram:az_wr_n
	wire  [15:0] mm_interconnect_0_sdram_s1_writedata;                          // mm_interconnect_0:sdram_s1_writedata -> sdram:az_data
	wire         mm_interconnect_0_epcs_epcs_control_port_chipselect;           // mm_interconnect_0:epcs_epcs_control_port_chipselect -> epcs:chipselect
	wire  [31:0] mm_interconnect_0_epcs_epcs_control_port_readdata;             // epcs:readdata -> mm_interconnect_0:epcs_epcs_control_port_readdata
	wire   [8:0] mm_interconnect_0_epcs_epcs_control_port_address;              // mm_interconnect_0:epcs_epcs_control_port_address -> epcs:address
	wire         mm_interconnect_0_epcs_epcs_control_port_read;                 // mm_interconnect_0:epcs_epcs_control_port_read -> epcs:read_n
	wire         mm_interconnect_0_epcs_epcs_control_port_write;                // mm_interconnect_0:epcs_epcs_control_port_write -> epcs:write_n
	wire  [31:0] mm_interconnect_0_epcs_epcs_control_port_writedata;            // mm_interconnect_0:epcs_epcs_control_port_writedata -> epcs:writedata
	wire  [31:0] mm_interconnect_0_cpu_jtag_debug_module_readdata;              // cpu:jtag_debug_module_readdata -> mm_interconnect_0:cpu_jtag_debug_module_readdata
	wire         mm_interconnect_0_cpu_jtag_debug_module_waitrequest;           // cpu:jtag_debug_module_waitrequest -> mm_interconnect_0:cpu_jtag_debug_module_waitrequest
	wire         mm_interconnect_0_cpu_jtag_debug_module_debugaccess;           // mm_interconnect_0:cpu_jtag_debug_module_debugaccess -> cpu:jtag_debug_module_debugaccess
	wire   [8:0] mm_interconnect_0_cpu_jtag_debug_module_address;               // mm_interconnect_0:cpu_jtag_debug_module_address -> cpu:jtag_debug_module_address
	wire         mm_interconnect_0_cpu_jtag_debug_module_read;                  // mm_interconnect_0:cpu_jtag_debug_module_read -> cpu:jtag_debug_module_read
	wire   [3:0] mm_interconnect_0_cpu_jtag_debug_module_byteenable;            // mm_interconnect_0:cpu_jtag_debug_module_byteenable -> cpu:jtag_debug_module_byteenable
	wire         mm_interconnect_0_cpu_jtag_debug_module_write;                 // mm_interconnect_0:cpu_jtag_debug_module_write -> cpu:jtag_debug_module_write
	wire  [31:0] mm_interconnect_0_cpu_jtag_debug_module_writedata;             // mm_interconnect_0:cpu_jtag_debug_module_writedata -> cpu:jtag_debug_module_writedata
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect;      // mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata;        // jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest;     // jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_address;         // mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;            // mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> jtag_uart:av_read_n
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;           // mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> jtag_uart:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata;       // mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	wire  [31:0] mm_interconnect_0_alt_vip_vfr_0_avalon_slave_readdata;         // alt_vip_vfr_0:slave_readdata -> mm_interconnect_0:alt_vip_vfr_0_avalon_slave_readdata
	wire   [4:0] mm_interconnect_0_alt_vip_vfr_0_avalon_slave_address;          // mm_interconnect_0:alt_vip_vfr_0_avalon_slave_address -> alt_vip_vfr_0:slave_address
	wire         mm_interconnect_0_alt_vip_vfr_0_avalon_slave_read;             // mm_interconnect_0:alt_vip_vfr_0_avalon_slave_read -> alt_vip_vfr_0:slave_read
	wire         mm_interconnect_0_alt_vip_vfr_0_avalon_slave_write;            // mm_interconnect_0:alt_vip_vfr_0_avalon_slave_write -> alt_vip_vfr_0:slave_write
	wire  [31:0] mm_interconnect_0_alt_vip_vfr_0_avalon_slave_writedata;        // mm_interconnect_0:alt_vip_vfr_0_avalon_slave_writedata -> alt_vip_vfr_0:slave_writedata
	wire  [31:0] mm_interconnect_0_sysid_control_slave_readdata;                // sysid:readdata -> mm_interconnect_0:sysid_control_slave_readdata
	wire   [0:0] mm_interconnect_0_sysid_control_slave_address;                 // mm_interconnect_0:sysid_control_slave_address -> sysid:address
	wire         mm_interconnect_0_f_engine_frac_cpu_chipselect;                // mm_interconnect_0:f_engine_frac_cpu_chipselect -> f_engine:frac_chipselect
	wire  [31:0] mm_interconnect_0_f_engine_frac_cpu_readdata;                  // f_engine:frac_readdata -> mm_interconnect_0:f_engine_frac_cpu_readdata
	wire   [1:0] mm_interconnect_0_f_engine_frac_cpu_address;                   // mm_interconnect_0:f_engine_frac_cpu_address -> f_engine:frac_address
	wire         mm_interconnect_0_f_engine_frac_cpu_write;                     // mm_interconnect_0:f_engine_frac_cpu_write -> f_engine:frac_write
	wire  [31:0] mm_interconnect_0_f_engine_frac_cpu_writedata;                 // mm_interconnect_0:f_engine_frac_cpu_writedata -> f_engine:frac_writedata
	wire         mm_interconnect_0_timer_0_s1_chipselect;                       // mm_interconnect_0:timer_0_s1_chipselect -> timer_0:chipselect
	wire  [15:0] mm_interconnect_0_timer_0_s1_readdata;                         // timer_0:readdata -> mm_interconnect_0:timer_0_s1_readdata
	wire   [2:0] mm_interconnect_0_timer_0_s1_address;                          // mm_interconnect_0:timer_0_s1_address -> timer_0:address
	wire         mm_interconnect_0_timer_0_s1_write;                            // mm_interconnect_0:timer_0_s1_write -> timer_0:write_n
	wire  [15:0] mm_interconnect_0_timer_0_s1_writedata;                        // mm_interconnect_0:timer_0_s1_writedata -> timer_0:writedata
	wire         mm_interconnect_0_pio_led_green_s1_chipselect;                 // mm_interconnect_0:pio_led_green_s1_chipselect -> pio_led_green:chipselect
	wire  [31:0] mm_interconnect_0_pio_led_green_s1_readdata;                   // pio_led_green:readdata -> mm_interconnect_0:pio_led_green_s1_readdata
	wire   [2:0] mm_interconnect_0_pio_led_green_s1_address;                    // mm_interconnect_0:pio_led_green_s1_address -> pio_led_green:address
	wire         mm_interconnect_0_pio_led_green_s1_write;                      // mm_interconnect_0:pio_led_green_s1_write -> pio_led_green:write_n
	wire  [31:0] mm_interconnect_0_pio_led_green_s1_writedata;                  // mm_interconnect_0:pio_led_green_s1_writedata -> pio_led_green:writedata
	wire  [31:0] mm_interconnect_0_pio_sw_s1_readdata;                          // pio_sw:readdata -> mm_interconnect_0:pio_sw_s1_readdata
	wire   [1:0] mm_interconnect_0_pio_sw_s1_address;                           // mm_interconnect_0:pio_sw_s1_address -> pio_sw:address
	wire  [31:0] mm_interconnect_0_touch_panel_busy_s1_readdata;                // touch_panel_busy:readdata -> mm_interconnect_0:touch_panel_busy_s1_readdata
	wire   [1:0] mm_interconnect_0_touch_panel_busy_s1_address;                 // mm_interconnect_0:touch_panel_busy_s1_address -> touch_panel_busy:address
	wire         mm_interconnect_0_touch_panel_penirq_n_s1_chipselect;          // mm_interconnect_0:touch_panel_penirq_n_s1_chipselect -> touch_panel_penirq_n:chipselect
	wire  [31:0] mm_interconnect_0_touch_panel_penirq_n_s1_readdata;            // touch_panel_penirq_n:readdata -> mm_interconnect_0:touch_panel_penirq_n_s1_readdata
	wire   [1:0] mm_interconnect_0_touch_panel_penirq_n_s1_address;             // mm_interconnect_0:touch_panel_penirq_n_s1_address -> touch_panel_penirq_n:address
	wire         mm_interconnect_0_touch_panel_penirq_n_s1_write;               // mm_interconnect_0:touch_panel_penirq_n_s1_write -> touch_panel_penirq_n:write_n
	wire  [31:0] mm_interconnect_0_touch_panel_penirq_n_s1_writedata;           // mm_interconnect_0:touch_panel_penirq_n_s1_writedata -> touch_panel_penirq_n:writedata
	wire  [31:0] mm_interconnect_0_boton_a_s1_readdata;                         // boton_a:readdata -> mm_interconnect_0:boton_a_s1_readdata
	wire   [1:0] mm_interconnect_0_boton_a_s1_address;                          // mm_interconnect_0:boton_a_s1_address -> boton_a:address
	wire  [31:0] mm_interconnect_0_boton_b_s1_readdata;                         // boton_b:readdata -> mm_interconnect_0:boton_b_s1_readdata
	wire   [1:0] mm_interconnect_0_boton_b_s1_address;                          // mm_interconnect_0:boton_b_s1_address -> boton_b:address
	wire  [31:0] mm_interconnect_0_boton_x_s1_readdata;                         // boton_x:readdata -> mm_interconnect_0:boton_x_s1_readdata
	wire   [1:0] mm_interconnect_0_boton_x_s1_address;                          // mm_interconnect_0:boton_x_s1_address -> boton_x:address
	wire  [31:0] mm_interconnect_0_boton_y_s1_readdata;                         // boton_y:readdata -> mm_interconnect_0:boton_y_s1_readdata
	wire   [1:0] mm_interconnect_0_boton_y_s1_address;                          // mm_interconnect_0:boton_y_s1_address -> boton_y:address
	wire  [31:0] mm_interconnect_0_boton_l_s1_readdata;                         // boton_l:readdata -> mm_interconnect_0:boton_l_s1_readdata
	wire   [1:0] mm_interconnect_0_boton_l_s1_address;                          // mm_interconnect_0:boton_l_s1_address -> boton_l:address
	wire  [31:0] mm_interconnect_0_boton_r_s1_readdata;                         // boton_r:readdata -> mm_interconnect_0:boton_r_s1_readdata
	wire   [1:0] mm_interconnect_0_boton_r_s1_address;                          // mm_interconnect_0:boton_r_s1_address -> boton_r:address
	wire  [31:0] mm_interconnect_0_boton_up_s1_readdata;                        // boton_up:readdata -> mm_interconnect_0:boton_up_s1_readdata
	wire   [1:0] mm_interconnect_0_boton_up_s1_address;                         // mm_interconnect_0:boton_up_s1_address -> boton_up:address
	wire  [31:0] mm_interconnect_0_boton_down_s1_readdata;                      // boton_down:readdata -> mm_interconnect_0:boton_down_s1_readdata
	wire   [1:0] mm_interconnect_0_boton_down_s1_address;                       // mm_interconnect_0:boton_down_s1_address -> boton_down:address
	wire  [31:0] mm_interconnect_0_boton_left_s1_readdata;                      // boton_left:readdata -> mm_interconnect_0:boton_left_s1_readdata
	wire   [1:0] mm_interconnect_0_boton_left_s1_address;                       // mm_interconnect_0:boton_left_s1_address -> boton_left:address
	wire  [31:0] mm_interconnect_0_boton_right_s1_readdata;                     // boton_right:readdata -> mm_interconnect_0:boton_right_s1_readdata
	wire   [1:0] mm_interconnect_0_boton_right_s1_address;                      // mm_interconnect_0:boton_right_s1_address -> boton_right:address
	wire  [31:0] mm_interconnect_0_analog1_x_s1_readdata;                       // analog1_x:readdata -> mm_interconnect_0:analog1_x_s1_readdata
	wire   [1:0] mm_interconnect_0_analog1_x_s1_address;                        // mm_interconnect_0:analog1_x_s1_address -> analog1_x:address
	wire  [31:0] mm_interconnect_0_analog1_y_s1_readdata;                       // analog1_y:readdata -> mm_interconnect_0:analog1_y_s1_readdata
	wire   [1:0] mm_interconnect_0_analog1_y_s1_address;                        // mm_interconnect_0:analog1_y_s1_address -> analog1_y:address
	wire  [31:0] mm_interconnect_0_analog2_x_s1_readdata;                       // analog2_x:readdata -> mm_interconnect_0:analog2_x_s1_readdata
	wire   [1:0] mm_interconnect_0_analog2_x_s1_address;                        // mm_interconnect_0:analog2_x_s1_address -> analog2_x:address
	wire  [31:0] mm_interconnect_0_analog2_y_s1_readdata;                       // analog2_y:readdata -> mm_interconnect_0:analog2_y_s1_readdata
	wire   [1:0] mm_interconnect_0_analog2_y_s1_address;                        // mm_interconnect_0:analog2_y_s1_address -> analog2_y:address
	wire         mm_interconnect_0_touch_panel_spi_spi_control_port_chipselect; // mm_interconnect_0:touch_panel_spi_spi_control_port_chipselect -> touch_panel_spi:spi_select
	wire  [15:0] mm_interconnect_0_touch_panel_spi_spi_control_port_readdata;   // touch_panel_spi:data_to_cpu -> mm_interconnect_0:touch_panel_spi_spi_control_port_readdata
	wire   [2:0] mm_interconnect_0_touch_panel_spi_spi_control_port_address;    // mm_interconnect_0:touch_panel_spi_spi_control_port_address -> touch_panel_spi:mem_addr
	wire         mm_interconnect_0_touch_panel_spi_spi_control_port_read;       // mm_interconnect_0:touch_panel_spi_spi_control_port_read -> touch_panel_spi:read_n
	wire         mm_interconnect_0_touch_panel_spi_spi_control_port_write;      // mm_interconnect_0:touch_panel_spi_spi_control_port_write -> touch_panel_spi:write_n
	wire  [15:0] mm_interconnect_0_touch_panel_spi_spi_control_port_writedata;  // mm_interconnect_0:touch_panel_spi_spi_control_port_writedata -> touch_panel_spi:data_from_cpu
	wire         irq_mapper_receiver0_irq;                                      // timer_0:irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                      // jtag_uart:av_irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver2_irq;                                      // touch_panel_spi:irq -> irq_mapper:receiver2_irq
	wire         irq_mapper_receiver3_irq;                                      // touch_panel_penirq_n:irq -> irq_mapper:receiver3_irq
	wire  [31:0] cpu_d_irq_irq;                                                 // irq_mapper:sender_irq -> cpu:d_irq
	wire         rst_controller_reset_out_reset;                                // rst_controller:reset_out -> [cpu:reset_n, epcs:reset_n, irq_mapper:reset, mm_interconnect_0:cpu_reset_n_reset_bridge_in_reset_reset, pio_led_green:reset_n, pio_sw:reset_n, rst_translator:in_reset, sdram:reset_n, sysid:reset_n, timer_0:reset_n]
	wire         rst_controller_reset_out_reset_req;                            // rst_controller:reset_req -> [cpu:reset_req, epcs:reset_req, rst_translator:reset_req_in]
	wire         cpu_jtag_debug_module_reset_reset;                             // cpu:jtag_debug_module_resetrequest -> rst_controller:reset_in1

	alt_vipitc131_IS2Vid #(
		.NUMBER_OF_COLOUR_PLANES       (3),
		.COLOUR_PLANES_ARE_IN_PARALLEL (1),
		.BPS                           (8),
		.INTERLACED                    (0),
		.H_ACTIVE_PIXELS               (800),
		.V_ACTIVE_LINES                (600),
		.ACCEPT_COLOURS_IN_SEQ         (0),
		.FIFO_DEPTH                    (800),
		.CLOCKS_ARE_SAME               (0),
		.USE_CONTROL                   (0),
		.NO_OF_MODES                   (1),
		.THRESHOLD                     (799),
		.STD_WIDTH                     (1),
		.GENERATE_SYNC                 (0),
		.USE_EMBEDDED_SYNCS            (0),
		.AP_LINE                       (0),
		.V_BLANK                       (0),
		.H_BLANK                       (0),
		.H_SYNC_LENGTH                 (128),
		.H_FRONT_PORCH                 (40),
		.H_BACK_PORCH                  (88),
		.V_SYNC_LENGTH                 (4),
		.V_FRONT_PORCH                 (1),
		.V_BACK_PORCH                  (23),
		.F_RISING_EDGE                 (0),
		.F_FALLING_EDGE                (0),
		.FIELD0_V_RISING_EDGE          (0),
		.FIELD0_V_BLANK                (0),
		.FIELD0_V_SYNC_LENGTH          (0),
		.FIELD0_V_FRONT_PORCH          (0),
		.FIELD0_V_BACK_PORCH           (0),
		.ANC_LINE                      (0),
		.FIELD0_ANC_LINE               (0)
	) alt_vip_itc_0 (
		.is_clk        (clk_clk),                                             //       is_clk_rst.clk
		.rst           (~reset_reset_n),                                      // is_clk_rst_reset.reset
		.is_data       (alt_vip_vfr_0_avalon_streaming_source_data),          //              din.data
		.is_valid      (alt_vip_vfr_0_avalon_streaming_source_valid),         //                 .valid
		.is_ready      (alt_vip_vfr_0_avalon_streaming_source_ready),         //                 .ready
		.is_sop        (alt_vip_vfr_0_avalon_streaming_source_startofpacket), //                 .startofpacket
		.is_eop        (alt_vip_vfr_0_avalon_streaming_source_endofpacket),   //                 .endofpacket
		.vid_clk       (alt_vip_itc_0_clocked_video_vid_clk),                 //    clocked_video.export
		.vid_data      (alt_vip_itc_0_clocked_video_vid_data),                //                 .export
		.underflow     (alt_vip_itc_0_clocked_video_underflow),               //                 .export
		.vid_datavalid (alt_vip_itc_0_clocked_video_vid_datavalid),           //                 .export
		.vid_v_sync    (alt_vip_itc_0_clocked_video_vid_v_sync),              //                 .export
		.vid_h_sync    (alt_vip_itc_0_clocked_video_vid_h_sync),              //                 .export
		.vid_f         (alt_vip_itc_0_clocked_video_vid_f),                   //                 .export
		.vid_h         (alt_vip_itc_0_clocked_video_vid_h),                   //                 .export
		.vid_v         (alt_vip_itc_0_clocked_video_vid_v)                    //                 .export
	);

	alt_vipvfr131_vfr #(
		.BITS_PER_PIXEL_PER_COLOR_PLANE (8),
		.NUMBER_OF_CHANNELS_IN_PARALLEL (3),
		.NUMBER_OF_CHANNELS_IN_SEQUENCE (1),
		.MAX_IMAGE_WIDTH                (800),
		.MAX_IMAGE_HEIGHT               (600),
		.MEM_PORT_WIDTH                 (32),
		.RMASTER_FIFO_DEPTH             (64),
		.RMASTER_BURST_TARGET           (32),
		.CLOCKS_ARE_SEPARATE            (0)
	) alt_vip_vfr_0 (
		.clock                (clk_clk),                                                //             clock_reset.clk
		.reset                (~reset_reset_n),                                         //       clock_reset_reset.reset
		.master_clock         (clk_clk),                                                //            clock_master.clk
		.master_reset         (~reset_reset_n),                                         //      clock_master_reset.reset
		.slave_address        (mm_interconnect_0_alt_vip_vfr_0_avalon_slave_address),   //            avalon_slave.address
		.slave_write          (mm_interconnect_0_alt_vip_vfr_0_avalon_slave_write),     //                        .write
		.slave_writedata      (mm_interconnect_0_alt_vip_vfr_0_avalon_slave_writedata), //                        .writedata
		.slave_read           (mm_interconnect_0_alt_vip_vfr_0_avalon_slave_read),      //                        .read
		.slave_readdata       (mm_interconnect_0_alt_vip_vfr_0_avalon_slave_readdata),  //                        .readdata
		.slave_irq            (),                                                       //        interrupt_sender.irq
		.dout_data            (alt_vip_vfr_0_avalon_streaming_source_data),             // avalon_streaming_source.data
		.dout_valid           (alt_vip_vfr_0_avalon_streaming_source_valid),            //                        .valid
		.dout_ready           (alt_vip_vfr_0_avalon_streaming_source_ready),            //                        .ready
		.dout_startofpacket   (alt_vip_vfr_0_avalon_streaming_source_startofpacket),    //                        .startofpacket
		.dout_endofpacket     (alt_vip_vfr_0_avalon_streaming_source_endofpacket),      //                        .endofpacket
		.master_address       (alt_vip_vfr_0_avalon_master_address),                    //           avalon_master.address
		.master_burstcount    (alt_vip_vfr_0_avalon_master_burstcount),                 //                        .burstcount
		.master_readdata      (alt_vip_vfr_0_avalon_master_readdata),                   //                        .readdata
		.master_read          (alt_vip_vfr_0_avalon_master_read),                       //                        .read
		.master_readdatavalid (alt_vip_vfr_0_avalon_master_readdatavalid),              //                        .readdatavalid
		.master_waitrequest   (alt_vip_vfr_0_avalon_master_waitrequest)                 //                        .waitrequest
	);

	system_analog1_x analog1_x (
		.clk      (clk_clk),                                 //                 clk.clk
		.reset_n  (reset_reset_n),                           //               reset.reset_n
		.address  (mm_interconnect_0_analog1_x_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_analog1_x_s1_readdata), //                    .readdata
		.in_port  (analog1_x_export)                         // external_connection.export
	);

	system_analog1_x analog1_y (
		.clk      (clk_clk),                                 //                 clk.clk
		.reset_n  (reset_reset_n),                           //               reset.reset_n
		.address  (mm_interconnect_0_analog1_y_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_analog1_y_s1_readdata), //                    .readdata
		.in_port  (analog1_y_export)                         // external_connection.export
	);

	system_analog1_x analog2_x (
		.clk      (clk_clk),                                 //                 clk.clk
		.reset_n  (reset_reset_n),                           //               reset.reset_n
		.address  (mm_interconnect_0_analog2_x_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_analog2_x_s1_readdata), //                    .readdata
		.in_port  (analog2_x_export)                         // external_connection.export
	);

	system_analog1_x analog2_y (
		.clk      (clk_clk),                                 //                 clk.clk
		.reset_n  (reset_reset_n),                           //               reset.reset_n
		.address  (mm_interconnect_0_analog2_y_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_analog2_y_s1_readdata), //                    .readdata
		.in_port  (analog2_y_export)                         // external_connection.export
	);

	system_boton_a boton_a (
		.clk      (clk_clk),                               //                 clk.clk
		.reset_n  (reset_reset_n),                         //               reset.reset_n
		.address  (mm_interconnect_0_boton_a_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_boton_a_s1_readdata), //                    .readdata
		.in_port  (boton_a_export)                         // external_connection.export
	);

	system_boton_a boton_b (
		.clk      (clk_clk),                               //                 clk.clk
		.reset_n  (reset_reset_n),                         //               reset.reset_n
		.address  (mm_interconnect_0_boton_b_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_boton_b_s1_readdata), //                    .readdata
		.in_port  (boton_b_export)                         // external_connection.export
	);

	system_boton_a boton_down (
		.clk      (clk_clk),                                  //                 clk.clk
		.reset_n  (reset_reset_n),                            //               reset.reset_n
		.address  (mm_interconnect_0_boton_down_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_boton_down_s1_readdata), //                    .readdata
		.in_port  (boton_down_export)                         // external_connection.export
	);

	system_boton_a boton_l (
		.clk      (clk_clk),                               //                 clk.clk
		.reset_n  (reset_reset_n),                         //               reset.reset_n
		.address  (mm_interconnect_0_boton_l_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_boton_l_s1_readdata), //                    .readdata
		.in_port  (boton_l_export)                         // external_connection.export
	);

	system_boton_a boton_left (
		.clk      (clk_clk),                                  //                 clk.clk
		.reset_n  (reset_reset_n),                            //               reset.reset_n
		.address  (mm_interconnect_0_boton_left_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_boton_left_s1_readdata), //                    .readdata
		.in_port  (boton_left_export)                         // external_connection.export
	);

	system_boton_a boton_r (
		.clk      (clk_clk),                               //                 clk.clk
		.reset_n  (reset_reset_n),                         //               reset.reset_n
		.address  (mm_interconnect_0_boton_r_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_boton_r_s1_readdata), //                    .readdata
		.in_port  (boton_r_export)                         // external_connection.export
	);

	system_boton_a boton_right (
		.clk      (clk_clk),                                   //                 clk.clk
		.reset_n  (reset_reset_n),                             //               reset.reset_n
		.address  (mm_interconnect_0_boton_right_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_boton_right_s1_readdata), //                    .readdata
		.in_port  (boton_right_export)                         // external_connection.export
	);

	system_boton_a boton_up (
		.clk      (clk_clk),                                //                 clk.clk
		.reset_n  (reset_reset_n),                          //               reset.reset_n
		.address  (mm_interconnect_0_boton_up_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_boton_up_s1_readdata), //                    .readdata
		.in_port  (boton_up_export)                         // external_connection.export
	);

	system_boton_a boton_x (
		.clk      (clk_clk),                               //                 clk.clk
		.reset_n  (reset_reset_n),                         //               reset.reset_n
		.address  (mm_interconnect_0_boton_x_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_boton_x_s1_readdata), //                    .readdata
		.in_port  (boton_x_export)                         // external_connection.export
	);

	system_boton_a boton_y (
		.clk      (clk_clk),                               //                 clk.clk
		.reset_n  (reset_reset_n),                         //               reset.reset_n
		.address  (mm_interconnect_0_boton_y_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_boton_y_s1_readdata), //                    .readdata
		.in_port  (boton_y_export)                         // external_connection.export
	);

	system_cpu cpu (
		.clk                                   (clk_clk),                                             //                       clk.clk
		.reset_n                               (~rst_controller_reset_out_reset),                     //                   reset_n.reset_n
		.reset_req                             (rst_controller_reset_out_reset_req),                  //                          .reset_req
		.d_address                             (cpu_data_master_address),                             //               data_master.address
		.d_byteenable                          (cpu_data_master_byteenable),                          //                          .byteenable
		.d_read                                (cpu_data_master_read),                                //                          .read
		.d_readdata                            (cpu_data_master_readdata),                            //                          .readdata
		.d_waitrequest                         (cpu_data_master_waitrequest),                         //                          .waitrequest
		.d_write                               (cpu_data_master_write),                               //                          .write
		.d_writedata                           (cpu_data_master_writedata),                           //                          .writedata
		.jtag_debug_module_debugaccess_to_roms (cpu_data_master_debugaccess),                         //                          .debugaccess
		.i_address                             (cpu_instruction_master_address),                      //        instruction_master.address
		.i_read                                (cpu_instruction_master_read),                         //                          .read
		.i_readdata                            (cpu_instruction_master_readdata),                     //                          .readdata
		.i_waitrequest                         (cpu_instruction_master_waitrequest),                  //                          .waitrequest
		.i_readdatavalid                       (cpu_instruction_master_readdatavalid),                //                          .readdatavalid
		.d_irq                                 (cpu_d_irq_irq),                                       //                     d_irq.irq
		.jtag_debug_module_resetrequest        (cpu_jtag_debug_module_reset_reset),                   //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (mm_interconnect_0_cpu_jtag_debug_module_address),     //         jtag_debug_module.address
		.jtag_debug_module_byteenable          (mm_interconnect_0_cpu_jtag_debug_module_byteenable),  //                          .byteenable
		.jtag_debug_module_debugaccess         (mm_interconnect_0_cpu_jtag_debug_module_debugaccess), //                          .debugaccess
		.jtag_debug_module_read                (mm_interconnect_0_cpu_jtag_debug_module_read),        //                          .read
		.jtag_debug_module_readdata            (mm_interconnect_0_cpu_jtag_debug_module_readdata),    //                          .readdata
		.jtag_debug_module_waitrequest         (mm_interconnect_0_cpu_jtag_debug_module_waitrequest), //                          .waitrequest
		.jtag_debug_module_write               (mm_interconnect_0_cpu_jtag_debug_module_write),       //                          .write
		.jtag_debug_module_writedata           (mm_interconnect_0_cpu_jtag_debug_module_writedata),   //                          .writedata
		.no_ci_readra                          ()                                                     // custom_instruction_master.readra
	);

	system_epcs epcs (
		.clk           (clk_clk),                                             //               clk.clk
		.reset_n       (~rst_controller_reset_out_reset),                     //             reset.reset_n
		.reset_req     (rst_controller_reset_out_reset_req),                  //                  .reset_req
		.address       (mm_interconnect_0_epcs_epcs_control_port_address),    // epcs_control_port.address
		.chipselect    (mm_interconnect_0_epcs_epcs_control_port_chipselect), //                  .chipselect
		.dataavailable (),                                                    //                  .dataavailable
		.endofpacket   (),                                                    //                  .endofpacket
		.read_n        (~mm_interconnect_0_epcs_epcs_control_port_read),      //                  .read_n
		.readdata      (mm_interconnect_0_epcs_epcs_control_port_readdata),   //                  .readdata
		.readyfordata  (),                                                    //                  .readyfordata
		.write_n       (~mm_interconnect_0_epcs_epcs_control_port_write),     //                  .write_n
		.writedata     (mm_interconnect_0_epcs_epcs_control_port_writedata),  //                  .writedata
		.irq           (),                                                    //               irq.irq
		.dclk          (epcs_dclk),                                           //          external.export
		.sce           (epcs_sce),                                            //                  .export
		.sdo           (epcs_sdo),                                            //                  .export
		.data0         (epcs_data0)                                           //                  .export
	);

	chu_avalon_frac f_engine (
		.clk             (clk_clk),                                        //       clock_reset.clk
		.reset           (~reset_reset_n),                                 // clock_reset_reset.reset
		.frac_address    (mm_interconnect_0_f_engine_frac_cpu_address),    //          frac_cpu.address
		.frac_chipselect (mm_interconnect_0_f_engine_frac_cpu_chipselect), //                  .chipselect
		.frac_write      (mm_interconnect_0_f_engine_frac_cpu_write),      //                  .write
		.frac_writedata  (mm_interconnect_0_f_engine_frac_cpu_writedata),  //                  .writedata
		.frac_readdata   (mm_interconnect_0_f_engine_frac_cpu_readdata)    //                  .readdata
	);

	system_jtag_uart jtag_uart (
		.clk            (clk_clk),                                                   //               clk.clk
		.rst_n          (reset_reset_n),                                             //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver1_irq)                                   //               irq.irq
	);

	system_pio_led_green pio_led_green (
		.clk        (clk_clk),                                       //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),               //               reset.reset_n
		.address    (mm_interconnect_0_pio_led_green_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pio_led_green_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pio_led_green_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pio_led_green_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pio_led_green_s1_readdata),   //                    .readdata
		.out_port   (pio_led_green_export)                           // external_connection.export
	);

	system_pio_sw pio_sw (
		.clk      (clk_clk),                              //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address  (mm_interconnect_0_pio_sw_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_pio_sw_s1_readdata), //                    .readdata
		.in_port  (pio_sw_export)                         // external_connection.export
	);

	system_sdram sdram (
		.clk            (clk_clk),                                  //   clk.clk
		.reset_n        (~rst_controller_reset_out_reset),          // reset.reset_n
		.az_addr        (mm_interconnect_0_sdram_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_sdram_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_sdram_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_sdram_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_sdram_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_sdram_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_sdram_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_sdram_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_sdram_s1_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_addr),                               //  wire.export
		.zs_ba          (sdram_ba),                                 //      .export
		.zs_cas_n       (sdram_cas_n),                              //      .export
		.zs_cke         (sdram_cke),                                //      .export
		.zs_cs_n        (sdram_cs_n),                               //      .export
		.zs_dq          (sdram_dq),                                 //      .export
		.zs_dqm         (sdram_dqm),                                //      .export
		.zs_ras_n       (sdram_ras_n),                              //      .export
		.zs_we_n        (sdram_we_n)                                //      .export
	);

	system_sysid sysid (
		.clock    (clk_clk),                                        //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_control_slave_address)   //              .address
	);

	system_timer_0 timer_0 (
		.clk        (clk_clk),                                 //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         // reset.reset_n
		.address    (mm_interconnect_0_timer_0_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_0_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_0_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_0_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_0_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver0_irq)                 //   irq.irq
	);

	system_boton_a touch_panel_busy (
		.clk      (clk_clk),                                        //                 clk.clk
		.reset_n  (reset_reset_n),                                  //               reset.reset_n
		.address  (mm_interconnect_0_touch_panel_busy_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_touch_panel_busy_s1_readdata), //                    .readdata
		.in_port  (touch_panel_busy_export)                         // external_connection.export
	);

	system_touch_panel_penirq_n touch_panel_penirq_n (
		.clk        (clk_clk),                                              //                 clk.clk
		.reset_n    (reset_reset_n),                                        //               reset.reset_n
		.address    (mm_interconnect_0_touch_panel_penirq_n_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_touch_panel_penirq_n_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_touch_panel_penirq_n_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_touch_panel_penirq_n_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_touch_panel_penirq_n_s1_readdata),   //                    .readdata
		.in_port    (touch_panel_penirq_n_export),                          // external_connection.export
		.irq        (irq_mapper_receiver3_irq)                              //                 irq.irq
	);

	system_touch_panel_spi touch_panel_spi (
		.clk           (clk_clk),                                                       //              clk.clk
		.reset_n       (reset_reset_n),                                                 //            reset.reset_n
		.data_from_cpu (mm_interconnect_0_touch_panel_spi_spi_control_port_writedata),  // spi_control_port.writedata
		.data_to_cpu   (mm_interconnect_0_touch_panel_spi_spi_control_port_readdata),   //                 .readdata
		.mem_addr      (mm_interconnect_0_touch_panel_spi_spi_control_port_address),    //                 .address
		.read_n        (~mm_interconnect_0_touch_panel_spi_spi_control_port_read),      //                 .read_n
		.spi_select    (mm_interconnect_0_touch_panel_spi_spi_control_port_chipselect), //                 .chipselect
		.write_n       (~mm_interconnect_0_touch_panel_spi_spi_control_port_write),     //                 .write_n
		.irq           (irq_mapper_receiver2_irq),                                      //              irq.irq
		.MISO          (touch_panel_spi_MISO),                                          //         external.export
		.MOSI          (touch_panel_spi_MOSI),                                          //                 .export
		.SCLK          (touch_panel_spi_SCLK),                                          //                 .export
		.SS_n          (touch_panel_spi_SS_n)                                           //                 .export
	);

	system_mm_interconnect_0 mm_interconnect_0 (
		.clk_sys_clk_clk                                              (clk_clk),                                                       //                                            clk_sys_clk.clk
		.alt_vip_vfr_0_clock_master_reset_reset_bridge_in_reset_reset (~reset_reset_n),                                                // alt_vip_vfr_0_clock_master_reset_reset_bridge_in_reset.reset
		.cpu_reset_n_reset_bridge_in_reset_reset                      (rst_controller_reset_out_reset),                                //                      cpu_reset_n_reset_bridge_in_reset.reset
		.alt_vip_vfr_0_avalon_master_address                          (alt_vip_vfr_0_avalon_master_address),                           //                            alt_vip_vfr_0_avalon_master.address
		.alt_vip_vfr_0_avalon_master_waitrequest                      (alt_vip_vfr_0_avalon_master_waitrequest),                       //                                                       .waitrequest
		.alt_vip_vfr_0_avalon_master_burstcount                       (alt_vip_vfr_0_avalon_master_burstcount),                        //                                                       .burstcount
		.alt_vip_vfr_0_avalon_master_read                             (alt_vip_vfr_0_avalon_master_read),                              //                                                       .read
		.alt_vip_vfr_0_avalon_master_readdata                         (alt_vip_vfr_0_avalon_master_readdata),                          //                                                       .readdata
		.alt_vip_vfr_0_avalon_master_readdatavalid                    (alt_vip_vfr_0_avalon_master_readdatavalid),                     //                                                       .readdatavalid
		.cpu_data_master_address                                      (cpu_data_master_address),                                       //                                        cpu_data_master.address
		.cpu_data_master_waitrequest                                  (cpu_data_master_waitrequest),                                   //                                                       .waitrequest
		.cpu_data_master_byteenable                                   (cpu_data_master_byteenable),                                    //                                                       .byteenable
		.cpu_data_master_read                                         (cpu_data_master_read),                                          //                                                       .read
		.cpu_data_master_readdata                                     (cpu_data_master_readdata),                                      //                                                       .readdata
		.cpu_data_master_write                                        (cpu_data_master_write),                                         //                                                       .write
		.cpu_data_master_writedata                                    (cpu_data_master_writedata),                                     //                                                       .writedata
		.cpu_data_master_debugaccess                                  (cpu_data_master_debugaccess),                                   //                                                       .debugaccess
		.cpu_instruction_master_address                               (cpu_instruction_master_address),                                //                                 cpu_instruction_master.address
		.cpu_instruction_master_waitrequest                           (cpu_instruction_master_waitrequest),                            //                                                       .waitrequest
		.cpu_instruction_master_read                                  (cpu_instruction_master_read),                                   //                                                       .read
		.cpu_instruction_master_readdata                              (cpu_instruction_master_readdata),                               //                                                       .readdata
		.cpu_instruction_master_readdatavalid                         (cpu_instruction_master_readdatavalid),                          //                                                       .readdatavalid
		.alt_vip_vfr_0_avalon_slave_address                           (mm_interconnect_0_alt_vip_vfr_0_avalon_slave_address),          //                             alt_vip_vfr_0_avalon_slave.address
		.alt_vip_vfr_0_avalon_slave_write                             (mm_interconnect_0_alt_vip_vfr_0_avalon_slave_write),            //                                                       .write
		.alt_vip_vfr_0_avalon_slave_read                              (mm_interconnect_0_alt_vip_vfr_0_avalon_slave_read),             //                                                       .read
		.alt_vip_vfr_0_avalon_slave_readdata                          (mm_interconnect_0_alt_vip_vfr_0_avalon_slave_readdata),         //                                                       .readdata
		.alt_vip_vfr_0_avalon_slave_writedata                         (mm_interconnect_0_alt_vip_vfr_0_avalon_slave_writedata),        //                                                       .writedata
		.analog1_x_s1_address                                         (mm_interconnect_0_analog1_x_s1_address),                        //                                           analog1_x_s1.address
		.analog1_x_s1_readdata                                        (mm_interconnect_0_analog1_x_s1_readdata),                       //                                                       .readdata
		.analog1_y_s1_address                                         (mm_interconnect_0_analog1_y_s1_address),                        //                                           analog1_y_s1.address
		.analog1_y_s1_readdata                                        (mm_interconnect_0_analog1_y_s1_readdata),                       //                                                       .readdata
		.analog2_x_s1_address                                         (mm_interconnect_0_analog2_x_s1_address),                        //                                           analog2_x_s1.address
		.analog2_x_s1_readdata                                        (mm_interconnect_0_analog2_x_s1_readdata),                       //                                                       .readdata
		.analog2_y_s1_address                                         (mm_interconnect_0_analog2_y_s1_address),                        //                                           analog2_y_s1.address
		.analog2_y_s1_readdata                                        (mm_interconnect_0_analog2_y_s1_readdata),                       //                                                       .readdata
		.boton_a_s1_address                                           (mm_interconnect_0_boton_a_s1_address),                          //                                             boton_a_s1.address
		.boton_a_s1_readdata                                          (mm_interconnect_0_boton_a_s1_readdata),                         //                                                       .readdata
		.boton_b_s1_address                                           (mm_interconnect_0_boton_b_s1_address),                          //                                             boton_b_s1.address
		.boton_b_s1_readdata                                          (mm_interconnect_0_boton_b_s1_readdata),                         //                                                       .readdata
		.boton_down_s1_address                                        (mm_interconnect_0_boton_down_s1_address),                       //                                          boton_down_s1.address
		.boton_down_s1_readdata                                       (mm_interconnect_0_boton_down_s1_readdata),                      //                                                       .readdata
		.boton_l_s1_address                                           (mm_interconnect_0_boton_l_s1_address),                          //                                             boton_l_s1.address
		.boton_l_s1_readdata                                          (mm_interconnect_0_boton_l_s1_readdata),                         //                                                       .readdata
		.boton_left_s1_address                                        (mm_interconnect_0_boton_left_s1_address),                       //                                          boton_left_s1.address
		.boton_left_s1_readdata                                       (mm_interconnect_0_boton_left_s1_readdata),                      //                                                       .readdata
		.boton_r_s1_address                                           (mm_interconnect_0_boton_r_s1_address),                          //                                             boton_r_s1.address
		.boton_r_s1_readdata                                          (mm_interconnect_0_boton_r_s1_readdata),                         //                                                       .readdata
		.boton_right_s1_address                                       (mm_interconnect_0_boton_right_s1_address),                      //                                         boton_right_s1.address
		.boton_right_s1_readdata                                      (mm_interconnect_0_boton_right_s1_readdata),                     //                                                       .readdata
		.boton_up_s1_address                                          (mm_interconnect_0_boton_up_s1_address),                         //                                            boton_up_s1.address
		.boton_up_s1_readdata                                         (mm_interconnect_0_boton_up_s1_readdata),                        //                                                       .readdata
		.boton_x_s1_address                                           (mm_interconnect_0_boton_x_s1_address),                          //                                             boton_x_s1.address
		.boton_x_s1_readdata                                          (mm_interconnect_0_boton_x_s1_readdata),                         //                                                       .readdata
		.boton_y_s1_address                                           (mm_interconnect_0_boton_y_s1_address),                          //                                             boton_y_s1.address
		.boton_y_s1_readdata                                          (mm_interconnect_0_boton_y_s1_readdata),                         //                                                       .readdata
		.cpu_jtag_debug_module_address                                (mm_interconnect_0_cpu_jtag_debug_module_address),               //                                  cpu_jtag_debug_module.address
		.cpu_jtag_debug_module_write                                  (mm_interconnect_0_cpu_jtag_debug_module_write),                 //                                                       .write
		.cpu_jtag_debug_module_read                                   (mm_interconnect_0_cpu_jtag_debug_module_read),                  //                                                       .read
		.cpu_jtag_debug_module_readdata                               (mm_interconnect_0_cpu_jtag_debug_module_readdata),              //                                                       .readdata
		.cpu_jtag_debug_module_writedata                              (mm_interconnect_0_cpu_jtag_debug_module_writedata),             //                                                       .writedata
		.cpu_jtag_debug_module_byteenable                             (mm_interconnect_0_cpu_jtag_debug_module_byteenable),            //                                                       .byteenable
		.cpu_jtag_debug_module_waitrequest                            (mm_interconnect_0_cpu_jtag_debug_module_waitrequest),           //                                                       .waitrequest
		.cpu_jtag_debug_module_debugaccess                            (mm_interconnect_0_cpu_jtag_debug_module_debugaccess),           //                                                       .debugaccess
		.epcs_epcs_control_port_address                               (mm_interconnect_0_epcs_epcs_control_port_address),              //                                 epcs_epcs_control_port.address
		.epcs_epcs_control_port_write                                 (mm_interconnect_0_epcs_epcs_control_port_write),                //                                                       .write
		.epcs_epcs_control_port_read                                  (mm_interconnect_0_epcs_epcs_control_port_read),                 //                                                       .read
		.epcs_epcs_control_port_readdata                              (mm_interconnect_0_epcs_epcs_control_port_readdata),             //                                                       .readdata
		.epcs_epcs_control_port_writedata                             (mm_interconnect_0_epcs_epcs_control_port_writedata),            //                                                       .writedata
		.epcs_epcs_control_port_chipselect                            (mm_interconnect_0_epcs_epcs_control_port_chipselect),           //                                                       .chipselect
		.f_engine_frac_cpu_address                                    (mm_interconnect_0_f_engine_frac_cpu_address),                   //                                      f_engine_frac_cpu.address
		.f_engine_frac_cpu_write                                      (mm_interconnect_0_f_engine_frac_cpu_write),                     //                                                       .write
		.f_engine_frac_cpu_readdata                                   (mm_interconnect_0_f_engine_frac_cpu_readdata),                  //                                                       .readdata
		.f_engine_frac_cpu_writedata                                  (mm_interconnect_0_f_engine_frac_cpu_writedata),                 //                                                       .writedata
		.f_engine_frac_cpu_chipselect                                 (mm_interconnect_0_f_engine_frac_cpu_chipselect),                //                                                       .chipselect
		.jtag_uart_avalon_jtag_slave_address                          (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),         //                            jtag_uart_avalon_jtag_slave.address
		.jtag_uart_avalon_jtag_slave_write                            (mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),           //                                                       .write
		.jtag_uart_avalon_jtag_slave_read                             (mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),            //                                                       .read
		.jtag_uart_avalon_jtag_slave_readdata                         (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),        //                                                       .readdata
		.jtag_uart_avalon_jtag_slave_writedata                        (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),       //                                                       .writedata
		.jtag_uart_avalon_jtag_slave_waitrequest                      (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest),     //                                                       .waitrequest
		.jtag_uart_avalon_jtag_slave_chipselect                       (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),      //                                                       .chipselect
		.pio_led_green_s1_address                                     (mm_interconnect_0_pio_led_green_s1_address),                    //                                       pio_led_green_s1.address
		.pio_led_green_s1_write                                       (mm_interconnect_0_pio_led_green_s1_write),                      //                                                       .write
		.pio_led_green_s1_readdata                                    (mm_interconnect_0_pio_led_green_s1_readdata),                   //                                                       .readdata
		.pio_led_green_s1_writedata                                   (mm_interconnect_0_pio_led_green_s1_writedata),                  //                                                       .writedata
		.pio_led_green_s1_chipselect                                  (mm_interconnect_0_pio_led_green_s1_chipselect),                 //                                                       .chipselect
		.pio_sw_s1_address                                            (mm_interconnect_0_pio_sw_s1_address),                           //                                              pio_sw_s1.address
		.pio_sw_s1_readdata                                           (mm_interconnect_0_pio_sw_s1_readdata),                          //                                                       .readdata
		.sdram_s1_address                                             (mm_interconnect_0_sdram_s1_address),                            //                                               sdram_s1.address
		.sdram_s1_write                                               (mm_interconnect_0_sdram_s1_write),                              //                                                       .write
		.sdram_s1_read                                                (mm_interconnect_0_sdram_s1_read),                               //                                                       .read
		.sdram_s1_readdata                                            (mm_interconnect_0_sdram_s1_readdata),                           //                                                       .readdata
		.sdram_s1_writedata                                           (mm_interconnect_0_sdram_s1_writedata),                          //                                                       .writedata
		.sdram_s1_byteenable                                          (mm_interconnect_0_sdram_s1_byteenable),                         //                                                       .byteenable
		.sdram_s1_readdatavalid                                       (mm_interconnect_0_sdram_s1_readdatavalid),                      //                                                       .readdatavalid
		.sdram_s1_waitrequest                                         (mm_interconnect_0_sdram_s1_waitrequest),                        //                                                       .waitrequest
		.sdram_s1_chipselect                                          (mm_interconnect_0_sdram_s1_chipselect),                         //                                                       .chipselect
		.sysid_control_slave_address                                  (mm_interconnect_0_sysid_control_slave_address),                 //                                    sysid_control_slave.address
		.sysid_control_slave_readdata                                 (mm_interconnect_0_sysid_control_slave_readdata),                //                                                       .readdata
		.timer_0_s1_address                                           (mm_interconnect_0_timer_0_s1_address),                          //                                             timer_0_s1.address
		.timer_0_s1_write                                             (mm_interconnect_0_timer_0_s1_write),                            //                                                       .write
		.timer_0_s1_readdata                                          (mm_interconnect_0_timer_0_s1_readdata),                         //                                                       .readdata
		.timer_0_s1_writedata                                         (mm_interconnect_0_timer_0_s1_writedata),                        //                                                       .writedata
		.timer_0_s1_chipselect                                        (mm_interconnect_0_timer_0_s1_chipselect),                       //                                                       .chipselect
		.touch_panel_busy_s1_address                                  (mm_interconnect_0_touch_panel_busy_s1_address),                 //                                    touch_panel_busy_s1.address
		.touch_panel_busy_s1_readdata                                 (mm_interconnect_0_touch_panel_busy_s1_readdata),                //                                                       .readdata
		.touch_panel_penirq_n_s1_address                              (mm_interconnect_0_touch_panel_penirq_n_s1_address),             //                                touch_panel_penirq_n_s1.address
		.touch_panel_penirq_n_s1_write                                (mm_interconnect_0_touch_panel_penirq_n_s1_write),               //                                                       .write
		.touch_panel_penirq_n_s1_readdata                             (mm_interconnect_0_touch_panel_penirq_n_s1_readdata),            //                                                       .readdata
		.touch_panel_penirq_n_s1_writedata                            (mm_interconnect_0_touch_panel_penirq_n_s1_writedata),           //                                                       .writedata
		.touch_panel_penirq_n_s1_chipselect                           (mm_interconnect_0_touch_panel_penirq_n_s1_chipselect),          //                                                       .chipselect
		.touch_panel_spi_spi_control_port_address                     (mm_interconnect_0_touch_panel_spi_spi_control_port_address),    //                       touch_panel_spi_spi_control_port.address
		.touch_panel_spi_spi_control_port_write                       (mm_interconnect_0_touch_panel_spi_spi_control_port_write),      //                                                       .write
		.touch_panel_spi_spi_control_port_read                        (mm_interconnect_0_touch_panel_spi_spi_control_port_read),       //                                                       .read
		.touch_panel_spi_spi_control_port_readdata                    (mm_interconnect_0_touch_panel_spi_spi_control_port_readdata),   //                                                       .readdata
		.touch_panel_spi_spi_control_port_writedata                   (mm_interconnect_0_touch_panel_spi_spi_control_port_writedata),  //                                                       .writedata
		.touch_panel_spi_spi_control_port_chipselect                  (mm_interconnect_0_touch_panel_spi_spi_control_port_chipselect)  //                                                       .chipselect
	);

	system_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),       // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),       // receiver3.irq
		.sender_irq    (cpu_d_irq_irq)                   //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.reset_in1      (cpu_jtag_debug_module_reset_reset),  // reset_in1.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
