��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%�����d^S$�0���<SG���0}�q�hS���.o�o�X{R�?9�x��ּ�@�����Y�v.'1t��>�1M=�\,�i�R5V[d���qh��+��j- �&u'h5��|�g����2\ǰɪr4Q����H[�Wlg�J+��1,Z��mX�Պ�$��0�s�zw�
h���4���.}�mA��,�d��e�%:�}�+��H������u����]�jז��S[�"Qc���qiS�kDj`��B�~j��P���"�͸Ii����=
{u�A<�x�f6�̫��BS�t@A�J%�ª�*�$L��d�3>��];��ʈ��$����!���EE��ђ�l� �L�#Lb���=���T�툠�1B��n+���&C�u�� >��"���;,�����7���3N��yr�>1�!��]���<?Sb>n�;��Ө��x��Sw�00n��B�a��:,�Ù ��!�۪�c�v2��n�*tC�>��<�.���U��rB���]��E臵* ʉ2 z�NQȲ#7��p���18���%�����Nk�c\�CB2�@5���:�tQ̬��G,�"q6x� n��C�A&�l+�2ަB��������1P���v
>U����a�q��b`Xާ��<�7�|��kA��f�<(� ǓL'���D��A�v����%�1LSmt%�����k� 5]�gQh���Ϩ�/ϝ9�)����{ٵ��LX�*�1@}��~�/*�1P|}�I�������LNtϹs� O����(E3�Pκ�_D�Y���=�����˛E�V��Xv
.���@�����P�7��(��^��&?��s��k�w[?I)w��L�$�L�|�mΌ�� 6�ƅ>�pL����]�E��ɇ�����T�Jf���~�Gn��Su�w�#Ҋ԰^b��"Ŀ�u4�DaJ�o��\A6����6/A��}n�f�X�6̗V�y%#�=Be^��[Cj�(�K3i�ݢ"�9�l$1=��(�<OldJ�jT=W����s�|7������/���z{�*�g���n�_�p����&�(�Hq�~P�<R������*y$
���]���G7V���+$8d��a5��Z%b�n5�P��SW��=3�[��h��*�rq����n�\I�[��)#M���7�?<�Y.�Z�Uw��I.���U��WіT8�٧��]m|e�r��� ��CN���	�i�n�Q��Fw������A'{ r�}�Ck iLS�Ϻ�+'���p�*%� ��+V�쩦 �B
�uI����s�͏<G�����\*�c�T
w;�p&���GZS�>��@ϒ���ݼ��ta{SޭM��Fj[�����_�X�ؾ�KW��9j(g�"�\����A��Cf��/�X �P�=�D;]mb���~%�� 70V��y��כ�-5/蘰��� P@׊m���d4�n�U�Î�7^����T���X�2Sz:,h��K��iDOC+&�_P���})9���$ӾB�o=��FS�dS{X�+��Ԧ�{~���-��"��{(��:y��&'�B�+=N�<Ǩ��,{M:G�=�lTK�� �.���l4�}Aއ�z�������g$���YU���_g��>��$uV��P�2���F+˔����L�t��l�O�����uP��#l%޹���i�����͉��ֆ��>�NDs�޲w�4�+�-��jM��0�R���>�v.�s7!F28A~i�#
61��>�CN�/ު�_�7��Nu�I�|��A �F���E����F�xYt�v!�@��*"?D�`g����F���{�ɜ1�m�$��,�- �q���&Y���������a=�?�zŔ�y�x;��q��k]2���z��S��ט��-vfLj��/?"��D5Њ>��A/��C�!eA�q@wkP&�ȺN�k�H����G��p��6q�jw)�ҩ�2�&�����/�?`��O���lφ}����O�'{�d�|�.��>ܕ�AE�����m�	/&��7�2�n.�d�*�Ŕq�%�n�����W��Zw?vv���m�.�G�̜<��qî7�ZǾ��T�QN��F�R��*����ܷ����˙�tG��6�����b)6��s��>a=���R�Fڸg�LnVb�
��e��@�̱+�Qxq���P@�8��f�8tynZ�����~��)�������ǐ�-�%>���p�c C w��qG���k�?�>��p]�hl����ԗ퇍B�}:�(GZ�3a�l>��0w����5XS��3�t�_j���۲���T��� ��m~�i.���8���|O{�+G�K*����0/\�\��Е��-��v��Cz7T�(���]�[��U��<نLv�<J�� �X �� (�ވ@��>��u;?{wz��A:B���Pt-7��O�?���Ų�Q������u%w���%,`�+W�p`G�%�*�]�G�&:)�9C�)��@*�j�q�Ͻ+��5ג+�Q,�\^(#i�B0,t�'�@E�DVQA�
��c�"�Ͽ�P��n��ô?�|���,�Mر�IQ xPz���O�����-"8�y�R���7����Λ	'W��]��^5�=i����P��: �\� �?v�(�I,[�ٝ]ޑ�\�g�u �Ksp�������5̒�/��
�Q�����X'�͒���ȭxWn����neBEC��MNtM�p�T��2��	vz"�@9T��8�G�2�L�ҟ�>��R'��V[��R=�h�G��J�>Y����n��LK�K�MX��N�w���n@%�X�]?Ԧc�:��r�bC�a�c���[���e���<I�	o���r�SD��8s8^XMc��<��EzHGz8�����梖���1�*�

>[?W�[uňa+�:s���	��+�S�u#�8�#}?�:-�g�$�Q0KR���y1���:��6,��=	 �4�Q�dC�����w�΅&f�\{��3�lrh�,d��ZVw!E��0NwԮ@{�),>F�\|��ˆ2%����*����)�@�;�t�!���ީ������)5Q�)��P�rZ��Q�N��F��y��5�{���������Q�"Kɹ�O�P�ht�Õ�'E�񛢄"���[�� �:*�Ho`�c��\�`xt;��x>�z��b�@e�U�'�y欕��_w8©���V���[h���ET�Jx���H:�p�Q��6���T�*�u"c���aaX8Y"t��f���C��B��v,|��ؖ��V�M�Q~�{�I$�N>��<��J!�i�_f��D8��\��M���I�;{^R�F�c\��,̦Á݁���������`~�sZF��1U�n	PP@����v�ٶ�WFmW���%e ݞWF���Z�C���X�z��{L�4AV4�'��zN�#�j��s�EzP���Z���F���G�#���ò�G|mg۸�CXe�'M�$M,��A�S�B�YQ���W[%�d���J�3MV�5�;�C�.����Ӛh��U�Y�Y���Ȁ������M=�rZT����"��0xQ>�M�4;vnJ%<���
Գ` ��Ԏ���3�̗@"紏���\����Lw���`�?9���lK^�1V��ȮW�Q���|{�Í�o��#�Mvt���4��6ᰦY��:>R$�ebA��M�g��ܙR�ĸr�H�����U��-�%�rA�����D�-�QMc\F'>ʰ(�_y�&E+{�>��dhfK�=D���b���v�AoM"ڼ���y*��R���F�(UR�v:@���(�:n�1$H�1kQ��%�5e���G�s�#bY5�;H~}�ڦ��	݅)V�E,j��`��嗊4<�������ĸ֣e��OkfX�s�P��۽ǣ;#)�����6�����
������"��1�)�V^��/Kj�hP�PKD�P�)&Y,��9#���d���qtpӧ���Ռ��T}�����GF�x������\��]�q%�bwH�v���6���-��#�w]�X'p���!���3ʥ�I���x��e�{���T����Qx<���S�Z]s�F{�%��˗����Y�)T+��kӭ*�DQU��$hJ��$p�׶��������7��A������i��'�r$T) Su��aL�=&�}�.��X�%(�8���HK����N��;*�b��{zw���&?��gXF\�����Х5�eKU7�O+	酦���l���<��i[�0@�D	� �jm����������sծ��~B�v�:kh�����{����)�nU����� ÈU�r�>Ky�����ׇ��I|�5�{<a\.�S�%�	�g[�#n�Wܕ*a|�����5������K��x���ףk
��|��3��G�F��g8�^JR��������/�X�
��*i�t�q�];��H��,�ߕ<V��)�F]P+�[�0�߻���:�d���t��g�m�:Nz�5�xW�u�����Ƚ1'�%,���_ڑȊ�zv��`���Ѭ�]2�����	�ߙƓ50�-4�fAF�/`u��"O��Q�o���"v�� BB�0�n��b��p�����Jзjb��>ؾ��)����`���,rH�F�x��Q�t?	��FͿ]�p���+��V�c!��k�\3u�L1�%t���ȼ��+�t�1d��W�} �ɣ�����=�֚�=f�N�����~�ޛ�P�tx�9pԹh���X�_�!P\@����k�T5��Ɲ�ln���o;f�b�e��ۨ����ٟT,> O\��L��w����@��՘s{�+�L-PTw܊�b^�?s����l�IZ{�RV�!5��GMz�brdt���랷���q��r��W]~ 瀢ڮ>���Ӆ������%��"(Hu��,�
���i�4�<�̦�6���iR"9����|h��Ư��f��GI�|E�p�ݎy�G���Ԓ���wh
}�����6Y"M@}@N��û���+�e"kX/d�ݛL�%v�#]��
���o
�\0� ��)�nU�ܬ�bH����7���I��3�}|�DBUl"�2l�}�z��S�$egK��ގ��4�H�߶�O�,��<��C��R�_�����x��
�+4g����;'$)Q�,oNGsu���.��0է��1
?�E��tɥ�s#��&ݦ�M�:f;��rP����P����"u��C?�}�y��A���7�{�꾐$:�t�CR�w^�����Ad3�B��$
ܰ'�e��O}N[�W(}_�����^���!�
�����Au�_V �b��Y���4�>���M׵F�A&۪���7]�(-����{BULOi�	�R�V��V߲�y�s�F8���tJĥ�H��F�3������W��ˢ�L ήG����ZOI+�ܮ+Π�OÛz`쒿���zh��O���!�e*d(ֳ������C�kZ�F���$��Gn�8�&��M9�A����E~��r��Cf�^"�Fnv��)R�~��Wn���2Hj���$%7[�t���:�����	������A���,zyԾ�V��m""ӳk��ς���z^�2��®b �7��l�oTvD^2ܑL��
� ~͵�z�{Rx���V�&���89�￵|/�[�lH�<��6��r�[�y�,d�_f��h�}��n�O����)d��c�����7]�t�a�׍FDx���(��Ꮿ�
��ݽ"�\gc�ֈ�N�coApCue{6a|B�$o�g�ܮa0�,���[��}(.���{���_|�m��,�@rv���z��Dɞ��5���v�A�c�!_Gc��H�:����Xڕ����FT�<J�p��{����{�e,�#(��_`(�Ocڙ�������J	�
�j����M��y���F�Q�)?����ja���=��1{�&������l�=(F�Щ�3��?}i�Z�|Y�)R�W)�1����ˎ�;�s~��ۛ����]~�a�2Wȇ��Y���x���T��bw����Uָ�$7�nW��<����~(A����=|٩ydݝ���~�[kMT�R�O��:���sF]�E����O�Y.3��_��c�n1�������(g��2-)Qd$Yk�4[ʣC�xl�����{�����+���޶ʿެ�k�шH$ ������*���
�
�퇡h���T�U�v:��&��Ŕzi�kT��ȁ�-��mpMB��aS�5�ـ�D�k�Y�b׾�`l�X���`�s>� jo-�H�Ċ=�4�!t�:�΁���Q^N�^[[�QD݁��z3`�8�����M8p/���z�5�z�<�L�P���h�W��$����٣������J��{�\��.�cu��d1�/sP!Q&��`��H����]�h�L}/���T��#��"�#���u����~���%.\?�x#Dw��2٥���S��� ��w=��Ң���0��p�ؒ� Rl������������KȂ�{�0��4�ĭbc,S(��У� �r�0�[R���R�`U��)�aJ[��"#?a��W�C����'��������)����>c^�A�UK7٪�ָ�X� 4�y��eU�.{�[r5.s�3��O0yF;���lq���DQ�.Oa�/B �`����g<�I���Lh������O��P���&WQ��K����
�H�mh�tn���i垎�^5�ul0sˬQ�"�r��}��U���A��Fmbydj��������tq)��� r��%in��l�*����.U��Z'�}�Cv`?����3��_��͍`:�8��2;x� �@��������S��aO������$�q��A��gl��qE�kt��vD?���X��cH&\~�6���f�r/�^�M�:������>_n�����ut�~R����fR��Ì���a,�2D���D�]�?��y��H �@�A�R��~�x� -1��*��ÿi���8����X�`ʵ�:N9�H�I��-��}RmR�c�Syq�^�����Ut~#��=aeZ�8��ūbK��i���������~��%fxxu� x���.A�UD0����.[�zTN5Y�G�e`h�ut����m)"�>�J�C���Ańpz}f��9��A�wǊ�)��Z,��]��Z�
R�Y����)�8b�o��n;��
i@�Ka�� ��x=����ل}l3�F{OdV4��<)W�:��3��T�A�2*'lD��5�'�]�e�[^ė������,~�(;��Zߋ8r/�5��	����J�{�g��C=��JrM]?_���Dq�pQ�>�R��zDw��9�d���3�қء�A�O1�l)x?���ܜ��IvA�9�6��16_Մ^I�z�^��hȤcr70iPz��%V*�n�ۗ�xˆj��%Xg- ��֖���)��{�3�,x�߸�e���4����b��5\h.�r2��m��)< ��Gp��%=�
�<��n3\���'_X�&.�R�ƙY�l+l��0�&eϖ��>��`�����^��	����S�c��6 �EX��|���Vl���e+I�="ڪD|��S)�O	Tmwl�chceV�Z�+�	Y��$�/BF��r���l#-��(��$]!��ag��U��s����FM�����wt<C�h�.���Pӱ�l�����u
j��p-�f�$��
c N�"M��(���Ϝ�T�5��-�vn��:E��{����*B :l��t�BR�-?�����47���@��Krw�+�g��m���n%/av1���,���3�-%ߦ�F�4���x?�mU�֮Ƴ"�8��M��
�&�5=�W�p�4��*@qѧ�c-�e��)��qI^m矎�4p.,��Q��r3/�c�a��߬\�9v����1�Y�����h���Q��5��01�8��2��6 fj�E}�qJc�#� @�`�Y'�<	�Ы�j�d�ȼ�C���J��)��o�q�/�|���7��L�&����C������?�����'�?V$���S���W5�r�=깬���}\zc��<���u���K.l��{M���z��K�y�W�����jX�@l��{�}�Cq,�߇^�6Nt�m��hچ^(��"K�5z�*�z$ìDA/Ev���bT^����ݎ�ېN�^�%p6d�l�D�����hA	"�e����#P��������d?P�/�ʭ�@x�ì����G��Ƨ��8�o��F�,Z�Z����P��ិ����g>h�%@��܌��\s�}�r�/����N4� �#ܬ�v��^.��L)nc�-%�]����]�0�$ˡ�f��DΣ��Bi'@����e���u�˃{��	i|�nqT�|I|����V�g��̧AK9�>�L�Z�N���cG$ɘ��r�|�ۯυ(�\��;3WM�K��a4�:��"���)���_�RB̖.�@�ޘ�`$�ri���(ba�F���N�D����l4<�ʲ���'��(0Ђ���08�iI�� f��2!�A����Y�G2�[��NX�L����Nݭ$V�:I%�!(skϐ�B1�����ʤç����D� ;t�,��
p�M���E�QE23ɝ��Z(����k�6�n�J��g���3�`���h���Y��H���r/V:u����p1D����P����NY�m C2��p ~�W�*S��h��(T�
-lx_>4�M�ph]����}���mP�',��ׁl�to	�>3��C�_'r>5�\�o�r:��+�D(���l\}��W�|m\��#�54:�=�@p�C3K�B�;�*pa\��A���4���^��~I���?-�y3Y��;m��Pɲ�_�*ݒp�(�6�"Z����%֖�r��V2~��@�� gV���Mks`2!��/\�Ƅ��N]�f_�k1�4�	�~<UW|)���$��/�7~����_���;��!g��*�
Y���){;��S&����E"�bB��)u?��g(�Vs)g�3��"Tw����U�!�]���u�Df�k��ݙ赒5o-p��0��*$@�q&�L��E�[J�M,<�� �M����REs|s%�sp��r?)c��8	A]Y��uɵ��j�u�I����se��� S�����F�Nr����[o�;:���0c�Qḑ�����o��ڽ��Q:��*�����gӟt��8���􎎀�`� �%���Ȍ�E�#�m��V�Gx��n��+������5�~fh���/��ə�G``��K�RD�	1<��J��D{VM��O���c/�#5���ۘPs��(�Ak1G�'J<edT��k'z� v�$6�ʀ��o���x�|�Y�}��?���~Z�G���ū�a4��88����H�l���t�m�ZN;�@8\�)���J#^m ռJ#���4������W[�Y,��e�;�Qc��
1��*���aAqz�D[�~
�M�0
�"Ņ�����7yL�&v+���K$|D �UE��,����ïO�h�8zhX�!P�I�`b�D�&$L��zxu]�H�<�w�����l�eBxY��+���m�Gg�}0�	#?e\�B�T��л��,tT���39�h��*�λG��o,�\��d�����\�'��+�G��c��W/�n�"I�"�Yq׃�,�J���!��{����g��C���rK7j�X[59���F���<�(����.���V�+$"!ھ��dO"�m��U���R�r��?P+��~��z]oC*��#�;���0��p�t��.��<��W�eX}�
e�чE��<7�ĳ��g�5��}Ė�6ʊ��ۯ,�E}�?�H�GE�ɋj��-PW���X�12�XF���"�D�0W��S >��Bާj���^�ƽ��-|Y�4��=�TR�}R�NdK�I 	�)�2I��-�s���8��Db˲q�i�ʻ�˳ӭaWa��Ѣ9���A�(��Ty�N�ip��ɤ����ڶ9>_��u��6W)-(6��*�.�Lz�&w�x����`<`��Xv�L�}�KH��]1�~�$�.y� ��V&+Et(T��BWLykb��8�!�i�0��A�ü���.����E �Lɖ��뫜W�M-��F��
9[�3~�3��|=�;Z�oZs��w#vR��a4��'͐h��E�&f��ܝ좔u�^S`�T�չ������ekQs��_	��|��e�5D�%�D�~5�k9���cV�Vz�*	1I�S�B�e7��R9,�aViz�G��m��&+�)3s�}�'�sp�M�r�V�'g����Nb�H;�#����x���(j��C��+K&���&wǠ� ba~��� G��� ��Kי��(tW-�j�o��W��`T
�Y�}��%�-�C��g�������a�P�O$�~cJa�V8n(�[Ƨ2����m���4�
�D��T���wp�v6̌ML5Z�'I��"A00���+���ގ]Ge�C�c���XɗL3�b�g�&�r@����FN�@\&s�_��)��q��BWx�����#c�й�Rp[k?B�Uvһ��6�»���^�����I�B�Y�Jf�P8��'� &�6ד>X��-��^�C5�@���D#��H��l<���s;�ŷ���5�h�"�'�g��Q$<�N)�?:O2@x{ |�G
�|x��� �g�DX24Yc��Q�]
x �0��ڇ���,g����lF�()����ޤ�����P����@�FhNj�!����f��4ݙ�D����$��D6S���1�ݚ�F��3�T��:�*a��e�Or(w���K��A�6h�ޮ�3;����]��i�[���"�
˥�LF�O���?�S���|Q���b,�f+kG�"��"�h���e�c~1_�
�؎:��A|ݪ�5i�BU�TO1���]��8-���I��>x:E�x�}K!�Tl8�p���w5qӺ9���>03H����q���fo�\0O�q��*r�N���rs5Im����	�;�>a"^��m����$�`Is)S��ޝ�W|�"���,n��8�`	K[�R/F�^�b�S��w��\ i/834�g���`�gd�:�vd�T�`��A!��SE����m��ኸ����g�y��	*��M����uZ�H�y:Íy��*�[��5��6�t������!l�7��:7���s\��PB��f���zR�$�49!v��H��/�osG����y���&�*�H��,���b�[-�w�Wep�7P}��#�fx9��V*B%��U��j~�N��Z��=�0z�$�I�)<���H�漆�����Au�"]�H�}G
��d��ǐ�.'9	�b��u	��w3�����~[/�I,iAY�[t.kc�si{AT�?�#g���{ǁ����U�y�i�G:��`��������Z��bwb�T�ӂ����:�nkS�LO���R���7�r7�)L��v�ͦ�zF��S0�B���4{y��ю��!��c�&}�O��$�-�ʑߌhZwz �'q`*�0�./�e��
(X4~|��Eh�b�S�ok+6ѶՈ�˘{�� �<~J�Wٹ���!T��╹��@�εL�d�*7�k�'dZ.i�)?ңA1�H�������b)���������.7\D�&�͔�x׍Nإzɓ��0���乀���]�����O����dٞ�VLŊ½V���� s�ۡ�'ʖ<w��&�1l>\n�p��R:2lU���B�h�+�+/�#�C#gB廃I����+5�t������_H���������q:�~�A�PH��x]��x��H��̚|B��6�y���m�/�@�����kg�����XMd�q�e�{���e{���v��Om?ym�jk�ȱ#~T\f��@�?n��(�� Z��QGzt�G&�fV��E
p�M矁K�s�`��B!=[�n)٦T�f��h���ː�-��k�hm7V��l+kL	 7'��G?b��Α��ly�����LІп�H����ɽ�ad�̴��?�O���5�Tz\����3�=3�ffkƆq�Vj���Z{�����ϻ�����99�puvWȰ�,�Ʈ���|Ci@czwl�g����$��}+�,�E|�s�����7ƞ�9������� ��@�D�Q�n��9�xm�ԃN�W��y��>w�-�y�|�G������dƉY7N��n!�N�<�9��>@�,�=��Rbg�>m.���[
e۽N��̟@��J��Ht�!����V�ew`���dn �%>�f�d6�b`m^���M��eg�y�&�'�����q����mu�(==���{���]B�4����B��Q|K��3<��T��/"�6GTZ'3�ɋTjk�ص�u�fw˩x����9)Y�]���KI��gԜ�&U,S�kmh2Ji�6�6��;�ĉ+�NӾ)��_�(�R��w������v��N9w���^ʳ 釿�/���7�FAWr�l���u3�Fg�Yu�(��enۋ��'cj\�C37 u_��9S��"�K�,�L ���$GF\�E���	tx�Q��پ(Nݺ<�)i)h�X�c`ȁ�Wu*��;��sv��bI�
vI�}㼚~Ӊ��x���LD��HTj�����ω�Y��=��N7�Ԩ-Qen�]fFA��@48<���N�������g<����k�FO���p:�U��i�k�d�dڙP> 왮����v�T�ꉵ��1BTޗ5��YZ�+?�/�r~���
�0\�T/,��2��T}>Ģ�d���zӠ;�2]��s��Yzo�Z88�qv�J��$.�S�~�r�J�� � 0��K����\�>�������e���]]�I��Z|�������g=rH���Ybh"�[_f��9u`9�l#� 5��L��nA2$=�_���;���C�&�+��_
����'�}4���z�V<�C�T\P��T���CD���29Ce+؆�_I�d����-��������=�@]�L��r�Xٔjm�{����W��Α��o�l 	�ވ��xh��&�W����m��U5�Pd|��n�]O|�L6���%q���b��v�:mN�&��yQ��)S�a04��X_���d�<�t>�:���q����m�G���_�/������g+��z3�e���,W�/�JU��#�=�<���2�c@>������2ٓ�8� "��"�F��,myX�H?�g[��\웯����e�X:�+��w���v�!0���Z�'/^���w�4(��gR�d��f��nq#4���.M�I���j����7U0�v?9�s��C;/!�����%����@>8�H�O�ǉ@dG�5)"�Ţ�~g;�mG�x��[�
9��*�ٛ�ay7)���
��şk��6h>���#�?��2��j��h��-3��#���(�r�Ue���CVdO���<�����ʓ�r{��&�������𐖄t�o��:3#Z�r�o���&kyU���x�����[b�=jΒ��C��V�^�ck���c�����ғS�X(�c�����Z�^�QB"fT_ģw�ϸt`���<�$\/�%���K��2M���%���J��q��9eu��q@4�X~���6�^X��k��$�˜��=�)�N�9įx�|12�Ff���t�#K]:��1�&K��-���xy9(�4k��h�C,'|�i�^��8-����&���n���!l��Faa�̂��-s�t���#����!�5�f�h�z:��~���ݣ .q� -�R�-;
�N�񹖿>}�(�2w�L��&+�.{ԑ��w몣Z.��c��|��M���Cb؀ER��{�(�w����5p9o�f�����V��Q0J�����y�w2����ӒE�K�*�V�!
�X��p�$'a��F��"���� �y푤�
��B��rN��J,�����C�H�aK���%j�˅�S��,X�*PS����_{��J�([m8�'ٯ��gv�����Z�[���u�&�hu\�><K��Oy}���?3�,�e0�Q*�YMǗ�R��>	�H�Qȏ�>��� �Qڙ�m1�Ƨ�������<��H3'kal�/����]�|�Pb1�
��))J~�����kl��/�f��ZI0�Q[�������q��h�ߺ�����'�"fH���7��]���=�4 gm��~��
x?�)�^/�!�� �B�ұ�cٯ���1��6C6A& ��苣�K��`_
�z(�ߌ���>X��ـ6�BR��B`T�t������iO4��
��Or}-=c�J��Z�j*��̏(�;q�m0.�7����$'�"l�ή���������`�'��d��~�ٛi�6몽���������7�'Qe���>��o:�����dk�`ٳL�-~Q�=���j���)-�IM��/Q��T@����DY ��Y��Z����x���`}٫�i_$PP�	���E`����t��=2v��/�fՋ���L�#M�(4�X�ÞjW-��OsX�Z�6���-8�1e)!a�eC�{��첎5wt0�H2J��ݔ���g���-^V�9Iħkǔ4��q���2��������߼kv��V���?�P�p+"cl�M0/3�����;tM��.9eҰqܐ��ʑ�C<�x$���0BS��b��@I)M��e��1[D��q�+Sh��I�.f�e���q�{C@n����� �=}f���q~$�X��jpn*���W��Еy>Di*�lO��'0�5�Ѧ�G��ٲ���"k������ٜ���j�4I��1(�t��'䖲�El�zc�����k�������T}>�â�$�p�Y�e(}�下�G��p�ϻ; k�:�]žUn��OoӸ�t1��0���SG��*K����$�0�̘��C���X� 8�yeЩ����G[��m��M��H%�R��b9KC��r��YR�PL���VQܫ}�̋9�ngmC�o�6n%W��+�8Əf�(om��
��:�li�He�g��������iM��adc�FGA1�]Kh�Cl;6����%j|�ch"�.{f��1��Lj�V\���G}��@|j'�?�Ss�}��{2�xw��)6���@����+b<2q١
�S��V}������$D��Vl�v��EvI?��P�Vy��#�[	B3@�Jy���捿���C��ER�)t"�F_x��k��zw�l��W��%����W�n�������gbf`��]��08�T��d���S�i�^��Q=�q%�76lx4\�1�B��R�+��;���B�	'lۥ䍻�J+B��,G���=�fKI����#�͔#ő����������(d�?�_�JG��V��]�E�B��m����S��i��Hۏ7�:v�#J8y$7ȭ���H��K8�z�~n$5���F�ܰ%����L�=��2�2>�m9i�p6�M�:LTK�L�q�I��"�v,[��Sv��Hx$��ȾcUk�<f?ļI��y�k�4�de��N�7�2�B�*;����h=���E~�:��%qh�C\X�~���*���������r����>���L*����%�'$���{n��=XU�x*��`���Oy�,�;���(�
q��9�b<����mk��a�d�Ь$P��O��;�2�ސIIⳎ�44�U��h�7p�f�������8�� [+�A&L�)�qg�'�p�\�BIF�_ex+=��.�����&9�q��z��e���Wj6��Bf�S�Z%82&7{�dz�*���5�p=o����\��"q�R��S:�zj4����IG6�mLv��k���,i����mE�1��o�W ���/�����.c���PJJBc��&�M7M�Iv���y�_v�o�r�Z�D�o����V�wK�ۧa���ƍ�M$�t�A܌��QF�O﹞D:�d"":�9�O�t�����"A�?_�@���w}zi�*����Vc����k*рq� s{�`�u��;Qž���Vx�B�-+���/�������5��x�k��9�m��%�o����C^�c'`ە?��͊ #�zᮢ��LK$������Nnғ*���Mc��w%&���d��eAp�!G'^�3k�[m�A�w�����BSB�i�R;�J����3��+l{����>"�����S}7�$d����P��!8`ګR��
9��cG&�1�����{+��������U��WU�;s^@�o��O<���t|=#ʈL̽q��
ţj{A�&���tm�U�8�K
\$l����MKW�"[���fMn�V�=+%������a���Z]a�ܛ��h���<�H%�TxR��Y+{6:��0b���I���ī&މe���p�9�����G�w�v^"L����v����ŞêeH�pJvo�ٵ��s��y&/�Wm�
{�%����e�P���FMD�*Y��2�S��]�6��w]�T��lq�,��d�a�f�f��`��s�2�UX� gx/���k��O¤7/g��bB=k��@�LG��}������T�%���_���'�Q��1�њG�v�b)n}��3�sF���e��������K�#�ǖ�E �ʶ2����L8j�@��j�c�Z��	�\�ߖn�J��2E�m��c��L��M�d;������{�,�\^����{~�& �f�S����"c��d��=q�3������\�=U���O���a#�(� �O;���T�������H���1��	�6gЂ�_b��6�����%�p��p��[8ڞ�`���S�9=�����g\&=����ϧDG�9��Kf�z$o�ޑ��8Y�DBIbҬ���?�O".G+�I�[��pe!{1IC�!/7�J_��ĺx ?��?�j<4���V�d �D!'
|�?t���9.��
{�W�:���栙^B8c�;����E��:}��O�P;��5�wJg�������K{�r���r)~���'��Ў��;٧��`�1�o��[�8���j�chZU��m}3F�zQ
�tgb_>4qQ�?�ɍdL������u�u"sU0 	�g�U5��A��x \�����7�]N��aٍ����
ɟ��=B�ґ����}���X/ZU1���� ��S�R�FuN���1]7D|`'=~#*Ի��B�f3�*��$kA�J�H�"R�d�����E��䣘$2r�u�h����	���P!�{2cO��o0�5�ށ��Udys1 }��5��F�\�[����)ӌRf���s���ˣ�|B����~�!9����;�w`�� US�,����0{P���#�:�Ƕ�;�}�TCc�d\�6����`
gt�@�����æ����v1l���GסB]� m~~�ں�8�DA�G�)z���&}Ҩ�[�1���I�*3eU��opX���YpH��nD�tA�	��5�-�$���DTa��pr�n�"7����|��=�QR�Hg;�R1�!�R�P��Zc~߸E��V+Z~yD��%M@q�|Ǧ�G{U�zv�χ��o�hϐ<�Fr�k��apsg2�y�;[����#�]O��]���=9�H�-����hc�Bu��m���f&��^�R	�.�j��P�k�wU���K�5�& �S��a	��tP����jq��gm�Q͇�4�^���7�w^|T�������� ԫ�&�5iw�: ��0�d�����4Y�f"Nxl�W.���h��	Wr��D�p#T\�wB/A0~V�d�� 9S���H��rʹf��}B�m͇��kzюE���Eѷ_(�����N	�
݅��U�S�����`]��)�z��첝y`!��+D�ߞ=*L�V�I�w���sz#29�T���'+#�R�MI���J,�o�E�d��7k��8��Yc�P�y_r�ʫ,��t��ɥ��,���>���d�;@�x������<8�Fi�Y�@vS\��҇�ia����Gzx4C�~D{_UO<���:��I�>���|��m�@��Hu�}��3ύ�H_��FL�f���4����s��N�>�FcA_uc�<��IТ�$��+K<Y�=��Ai$��)���*L�OF�ܑ��Rr���΋��'�s51��o���-B��s_����>�I�҆Q���P��G�����u�0��42��)�}�J��~-�3i^��|��3��SA��2b`O۽������%���V��nc�vƉ�7�8�s�-p�p?��EX�`3A��5/�dðz�1���Y��w��<L���-�ȘIJ�s"�mҒ�}Ԙ,�]�6gvR�L;�xM|�
������*�)��9��F�`H�+�!��@���Y�MԧY(��y�u�MmҀ��l�d}��U>��]]ܔ�(�Cg̍@l�1����cU*��ۛY#�s5�����ib�h�g��QӺi���S}Nw��[�4�:�M�@
����ഥ�@?"��E��`28cѠ���"Җt��%���)#6ܕ���1����6�>�XVZ��Z7����K#����|!�i~�Tq?�ʨ��gK�����>l80��4"2jl�$O&+{Qx�$��Z�_��2��;�.�Z�9Y�>|O i'��T_5@�/��7%:I��[�t�g�����S,��/��$��?{�!�|}�t
X"$1%+�S��WQ���[�<���6=��K�}�i__�竑X�t�
]�_�3@�0>�	'�l�ϧ<��W����〽�?��])�o&IT�-sӘ}�>}�g�f�����שn��*��D������r����'pkDz�g���!qe���T�]^_,�qʱ���?m�Ό��g<a���؇
xK�_FrQެ=�LmP�9���%<�	�n��(:
��'�������[�Fq�� ���ƿ���'�V
�-�g�h�0�r�M1��k4i{Uef���m�E�*u<s.m��*�u�D�������a�}�������/q���w��֚����UE�X�r^�|l����"*�9�*X��B�,�6u�����xsM91o��}o��|�#8>�m":r�n��?� )���lv���ݵ�Z��YV��[�ƭXz�ޮ#��m��'�z��$�k��oj�����ڦ-�~EF��M�:+�(O~�+����{UŠ��}ꩡ�A(��v0�X��)n
���^�������S܆���{w�&l!��*O��"������u�l��5EE�L���c�T���)<��w�$���@��s�Ԧu=E,�F�W/����Ӕ&�V��n���	I'������[Y7�XL3.^/���Jqi� �#?�ݪ^ĕU�	"��w�֍<l�^��5$�Y3XX2��25���oP��"�����iWur����wV���p�RG86��yH��|�5�4�����zd>��tpC�sp��%���3�J�)����!Kw2H2�~��*p^p�c_!�j�;Й5� �0�9�@.0�+Kާ�\��i�	؂�D�F(�`��"!�������Q�~��4<���OM!���������u A��������8hwfS�Kb_�f� �����6��9Γ���7��Hc��<|!&�����L\��x�:��ga����/�@E�_��K�RY�i,'�x��c~�z�^�����	l�a0pΘ-� T��
ԽJ��H%��l	G���j�>�O���Z�̉{���&���UoF3P �<gt�F�
5�� YCBlV~xJ���H6��J����ѻ}�/P9DbDoR���άh��Ex��ٵp��0��'��C e_Wz�v&t�:8�W] d����(5��ñ��j�����3��.(ڲ�ɮrs��c���ݲ��7.�`�!�~�y��N{��X�6�A��L/��� �4����I�a��j��/����߶&B��Fn���&;�qD����{�߮�R����
�8;�S�1k�*���(:q���?�r2�oS	ueSQ�R���ugja�i�%`Ӥ���U�ţ-;�j/�h}~9��fr���g��1B��^}��<���:�s>�f8R3�����a�i��zN���Vg�k�o�Q�#�<j�<��"����Z�+m��ۯ��(�"\��q^�mʦ�7��]����ȷt���^d=��$_�l4S��2�س��LE��-�jNh���:n[i����	�&���o�7�H��7g)��l�>%?)��N^$��h)HEϧI�_9�MN��n=���(���\M>�A�~�RB�c?D��K��RSI����@B,�T�Sy�<Z�L�*;��-êe
�q�*1�\0R0V���$�������I*�.V6w���S���ή<r����H�%7֞�\����[
?�E��IthP�ҙs�	J,pi{f0�7j�Q�h]�B���Y�����ӈФ�c4M���$x�F�c�Ze�95��P��HN���Bo	�:_�Նr��\�H}��5+�Rh�d�)\Ek��L�|�p������A�F
]��dKQ�ޞ����ԃ�P���~dfcڎ+O�6:�)�T�ˌ���{Y��K棯wEr���gψb��JTx�-{�dm]�:`b_�8×�@�5�����i��ɬ���qO��%�n��E�����`��o��S��ű�>�PV(pX�t���2��r��yͨ�K�������\(�%��S%�F5 �����f�v��.׳kS���9��d�����Hh8��Ow�i%���<����z���R�;.Y���7�9��	R��@��:BA��W/PFd�g��S)�u�h*�	nQ7�^yx��f�q��` ����fRl��g���JA�C��[}µ����g{��E:N�݁P����l.��bث�L�l������1Ius��J��(���|Q�5�"�sԭ�f������he&�%�1e)ê��m�%�����yN�|��^��cbU��\���0����zSw)�T�氥�7)p��>T��rE��a�f��X:6�6���|e�4�L��P�}I��D4l7�sм�����B׹SR2J���s/���&�,�
*K��F�70/�;cY^���F���;=k�����9mْ(�i���l�#����x��
������7֯8ߪ����.J�.�'V�a9 R�X 䈎��8��bAw .򦋺�bc�m���tSS9nr�ʋ��v��#0bJ�TV����hB�����O�~ZM��r�2!����}$0 ڴpTnG�L%���{��a���!' �&c;��dt��كF�����.ky�p�*�Qº��'��z�:�9D������A ����Z�������ݵ�C���S�fS2>��[�ӷ���J��G#����g��z����������kğ+/��,��ܶМc�Y���}p���^���7b�#�N�7��?�]��z����0Ai��y���x%��kV[>�K����1ǔL� 
k)N¿�:�;�9qM�_{�ӓ\�?��~�d�A�d�RP%���$�V����7�V�}8Ѽ���"ޜ�}p��U�c��A'\�R4���S�	=9_��?��á�+#��U��`������~;&@��dp>(p��> ��)F��[Kġ6S�R������J����*x�a9�3ar�2I��c�ny�D��N�5�y�����/�=� ��硎��&½-w���:"0���D𾆼�/�3�!�x~�� D/�
��Dw�KZ��+wSo5��\<㧜\��?��?U�_�0,�Z'+]�5�ei��9�E�!�`G
Y�c|-�5��������\�9l��� ����'\�K�B0���^ƣ�y��t�%l�;�.��j�9�	���Jq�����(���|��?"�}6�I��Xz"�y����'�R��U��GT�T`��*ihjMP�xǊ��i��U�j��~��?���$��A��|��)�p�Z-�9�vZw�-�KB�8���0d�q��;���^��)��bw���P8�����j4��␔V�J%]E��~��p�d���(�Oh�5'P.���:cp�y~�7�f�o��tY�*_g��&�.;�㔠��D
>���Ǭ?u(9���&��n�wp.ttQ�l�_-�UC��W���ĲZ�#����"����9e�������-H�p:�ZP��:a@�~�D�m=^�
�J��0-�Q���5h;��@N*B���E�<X'�������4�4��Yl�s]_J������K<��������"'�;�"����O�اZ�0����&������=7���jFK�Ű�
o�m����m8��q9�pi�G��>���XN/��멼��zFU��<ޓ�9��Bd����珫�����u�w+y��X��kZ��?��|�մ8�u_f����Ka��=��3}L�dv�DT��Mn���mȀ�"�G���f�ؚ���H��0�1V�mwWa#����y��tͦ�fqB����3iTr�J*n�r�&����:S�UI�X�2:��,��
�9q�<�AN�4����}]�8���11��t�;䦥I�_%����V!@���5��&h�Q�bV2�C�X=P'��]W~h������l~��4�_��]8t�d���wPqj���4ouX
`��� �^��ja��0rw�'m(h��4a9>�[��=�$�_V����k�~�5�'S�fi��Ά�����eb�]��B��"��YQ0]{zD���>,���&������M����4�W+��f�i��	�D�K�6YJ?n�6�X� o&��<�օ=$W?�_͋�9[���s��o�ptc��Я��H��_���&x�դa���S�O��V#����0�,�ѩ�2�oմcy�H� �D�t�gW ��ơ9W�c)уtB>�5��o��>��NL���V��r�!�h:�px�Lׄ�*U�E#��r�7�w�������TR�d���Q��[��>�49�f��!ݴc�t��A�����x+�[c��sxrbY0��O�99�xU�GFT[jrq ��[@��)�����&2K�8��`lY�M~f[��M�,��?�B��X}�N�J�G_ø^B%:j����;�9=XŸP�hN��i��x�1��A]�"��yPP�T��MOG�^��NR��V���[,��o�.O���P�C.J���2,��X���8F���'kv��/�E���A��R�G�e�{/X*n^\f�Nz��:�"�I�.50���8Z:.辁�����{�(
?M+<Ϳ�ͺόAl�c�
t8��G�`@Vʰ�ci�¿d�͝�McQ�����8�yl��pАՉ���@	�u`���G�8伺���9��_ �tI�9�Z�5x��F(�,�3.�zvI`��a�g&%b.���xb�� yq��,�UіQ���A����5�
��X���xҐ���ꇔ�8��=A��k��ʏ���ЙO5'�k���:ڀX����5���wQ ��?��jŠj���&�v>/��a��<�4��ic��w���3��6��	��A�[��4`����w��ws����CI�$Eo��6m�i����bZD�O��P~��wR3�zG�����[#�s���#��K\��z��=-T��;����n�To �p�G)g��;�(�#A�TEMm�� 5e`�t��W�r�%D�uh�Tbe�bn�Y����e�:#_��(�4�׍ϯ��ꥒ<�(�-�|�{$S�;`O��9p��{<�,��g:{N�}�������m4B��:1�/Zr��T�~AM&k��_u����W8�g��\����;��A��n��J�Y2yO�R2��꣟f�KU�y��@�r$	�1���7�t'�H�ٽ�['�s��~̵��M�'z=:��l3oK��
�B��v�E?�����}�U�G��۱�����%�%�+����.�FW�
��@t_-�گ&�ސb=�T!+���|l�e��0y�4�]����E���ME8�=-+66(̸k��:��mP��7.�o�j��?�@�V"�T�=��j�(�����3xpV%]@b���q�e�!AE������E�M�-U�І��L Ks'�٠��%3�`Q!��n �����`�
�0=vG�ZZԠ�r6��!r��d��Гm|�f���?"��MJ-g��O��9vVr���N������}^ܔk೎X�M'���X��!�޽��B᠜�+&d7
�b���O8Qq�Q�5�8��������l����Z�sR1���55�{�>̖^{'��@B��O�㲕HY]�{�#�T�L�@�^��!(0����g��^��A�5���;�޼-ߢ:쒼ȉB�C�����]8|����z�#�S\:�;�п]�.�I`^։�hL9��2�r퓍b�p����K�hC_�Pv��R�Ͷ9��O��?I�)rD����|0�KgQ��M��e��d��`i���7w}���Hϝ�5���4(��'���󬅀N��;���1�\���������<�=�� b�J#�(D�.g�#�%���Lr}�4s�#`�p~����,��S�A�$ ڱ��;�H/X/�_G\�s^C�r�3���\�E(C�0��&h�2��_�������`��6�xa�Y$��ƃ).��m��:�f壂��g���7��P��#*�~q5��{蓳�#'�
5\�v��ڏm������	��o�����6'ۧ�oW���r�I�yzֻ�ǉQ�(��rp�v�Z3�gb��Ef���� ��m�q/��f����L
�x*�Жog���Ԋ��/��GI�����݊�?W��!��$D��	16?+�f�-E��oɞls��X>�w�r?<hT��b�}�' K~T�	mg3��Wc�U���������h8������D�u&��Idg�I�n�{X��p�Dc����f�=
n���7��`��|\67�g,Z��(c&��W����j��5`��j�����llr��P�E�E��O��+ �O�Z'��m[��G�z���PH�;�(C��fo��2	���]e��'\aFTw�����Ys�A�t��<�UN���)1tQlw���m�����7�d��7��L�`1�68��ޢ3�Ĝ�W�,�ʘG���[������r}z�Py��F��Y��������!&�g�'���y�lj��e+"}���N옱$ �Rڕ7N��IG���csB�����#���.��f�h�`@��չ�_֞+�3]h��Rkukb��х�YP��5���B����>F�٭��r��3$�E�Ea(��:;_w�{����V�l���(,�����rtsآ�ݒ��Y	)����A�s1w��D���"l���*��g�8LH�R�ǽ���XB�U�迍،��l���}5������ػ���7dS�������K;����r�I��=��%j����!\�{����#~�L�-c�'�2�V_�Cd���g��h�����x���Gt�yߌWX�����̚�oQeF�iPK;�h�$)8�J�bNT�M�4nm��w�Ơ�C�Q�Տ
�`���l�g�/�7��~B]������5�f��ԍ	b� �����[Sr�\�V�)�2�k�c�΢2�WH�6�1M"�5?:lᡁ����CS
����S�yx1Mjx?X:n6I�q?�A��b�c�Y�»�Iz���wvk#�mD����([��!Mwk/��z���D�ڷ*v{p%Z������ ?	>��r,���:��@�Fe,��\��x��P�pD�A��Y��47eX�!)�v��Njl��N���HބqRT��	.����xy�[���z-��}�C��ݶ��iď�̪ż}r��E� �1��]�[�E�L�̃pOVȏ��0��]���lCvU��eQ��e4Knԡv�tT��Xd�!��2Ԥ���VݛzuŉPf��+���yޟ��Ԕ��,F�.�����Lj;-���B|ƶxZ�)��C��e�!#>Ȏ�p,ԫ��!f�N����\�	�3�����~Ihg�ŷ��QAǸ����̘�H1z�&ϼ(���T:��G��nW{�r+G r�iR ,��I+���K5���hR,�zEqAY�Uɩ�`��R
BY��|��3'��D MD���o��)�7!�R�ŁS��]����I���ye7;?t:�r�x��(�ş0�����������9;ccˠ0Ŀ�`�C���y��1T����B���杣*N7�O�_=��3�1˅ W�B�=x��w��1^{�৘F�Ø�Hl
P������L���n�V�Q�D� Q� [��z'�t��ǩ�����{��uK�V�!Ӣ,� ?4u\P ,���|�Li�C*m!l����"�6Ֆ��>��"�N�W�̈́2�V������̘����ܠwF'��6�
+��Ɖ�C��Fw���'����y�N^3��c�	j�c-za�k�=�t��2�C:��C۽�e�(���0L/�r��Ȣ�4گ�:w�����g1_Ǿ�s��`�b�Yo=�;}�j��R��'X�IS>�W<��k�ѯFG��a�m1��5S��9�3���csM���
"��FF���1Mn�T�R�Ji��	���k�41�p-�|&�e�j���+��+�Nc���s���f��X��NS��,�P��!tE��.^��|�N��(�L8�Mձ��U:Ev��Gh�i�Yv4��KK���M�/D�m�͵/�e���U��U�~v)4^[k)�gz������O�?��s�,��s�"]�������
��Ʉ+��A�hJ��>>e[�l(lt9��ͣ0\,�.��Ύ��9vގ���<i00�+�ˇ��JB��nGv�9�yM��p͈�'S�2��.�N�z�B��&�d��OO+?�Db�I=)�j\8��?x8kB��Ev-� �^��K�婑�q��yW"W�>���c������� m_
���=��÷�f� k;������yGg3�[S�>˜�шJh �p��@Q����� X��ٷ��H�W���&�r�[���u �L�jiĩ-A3P�Y���q:���F^���i	���m�ėq5���6��V���Ʌ!�7Ʈ��������!s/)�����R=�:�Z.&ALQ��[Д�PP9�z}����@ue:�ӻ$F�ު�X��@�r��t����$-\��9b�KK>8�D����8"�g��0597��T�r7��^��L��
0�FlR0d��im�L�,Z�_�L*~m�xl3dmp�8�>D�]�C�*y�p�jQ��z��f
R��.D��݈�����]�mT����i��Ap�����G͊�9�fiS�)|RN(71�{��a��Bv�.��*�� �,I�$ֈ��>5�A%���a��$]���n��-B�����ڢ��퉃�t���۾Y"8�{��u��5���E����KƆe�\S�DUAmy�Ωg�]���P��U�F~�k�(�v�#5SVR�$�j�
��G��t���a���8�����"	&���1���o�Ќ�TL0�L����#gzk��sS�x�W55���,���δ�=�v�D��K��Ɵ�q�M���WvaVȱ�@�
d�,������S�G7�lT�?D�yW�;.�Ԉ�k�o��t<�p��i]�K�x�Wj8A�Dd�߅k�H����`�}%�>�j\i K�_�ա����3� �;^�mN ;�u���^iZɫ�EGJW��+ꝍZ�0��o��?� ��
��(dSR~dPkx}:�W�;�h�Ƃ
�e�.������R�&��Lu����D8����O��^=�o_�7�g�� SaD��qZ�o��&��]�bY���,�I�]�zcgK��r5|,q�sy��,?vt����Ib��r�ǐ|����شn�����G^�	����6/5t�*��.���_�CCʧl�-�p6.�c���yW���8�v�h��
��Ѱ�I�PBI��.Ñ\��
�>q�i��cb�^�P���g`���		{��4֐�����*���2����6w�8��}W�}sȣ��J�dMd���dYw(��2��{�\�1}_;�Ӂ(�4}	�%dzWW7Y��z:�\O�/v��/h�_��wH�p���'��j�a��F~�@tJ�"�j��������ؾԚOx@�������H}��R�j��4�5`�ƞ��Ec@C?c�h!��pJWw0��@$Ek+z{�?�4�&�k=qt-�BRۀK��Y!)�4��/c��$VU�Ud�?��� ���Ć���
�n���6�D��;�ΐ~��| L(/��
�.�M��b{w��I�j�F�g�At5�_��oH��&ti�D�ܥď���U�Ԕ�|e�X��h:�w>%��=�`�������E*����s�~VTk������$�d�4f���F7�㘩	�W��`1	`�{PNP
w�D3w��l���%����hq����6��W�<��t�T�8-))Cb�!��Ոs���Vrk� r���n�Q�/j��N<�+���ʥG����Α��B���ߺ^��
{���T;�MW�K�GB����um��g����h��}�+�q�r'WqB��K(�OC��Gk�k��Y|�'b���z��T���8 T,0!p���}�jk������K�ƚ"$�5�
ձ&�M�y�x�<��O�/�C_��RN=[Л�(�] ($�d��l�A��r�._��&<m��I]����!!V't���^�����@�M��������;5 ����.�)�g��b�׵��F<ө[H�Uq���
�\��2R�Et��C�\�?��SQ�xn՜��ᵀg��g�Ee䇃��	m�\�So'�Q@#�W&T{9��՗�D�����]����w��9�LH�HTX�-p-�����V�e�U53�w����z���Q��<��7��>�������$W=3�-Zk_>We_EJ�5���A=�6u+��D9@Eg���`M��ih6�N�)c����.>�ef�.���[��n��2=�4c�}���y(���ނ�&�V���Q�M�,�^ �����!ᾔt͋�6���r�8G8rNy�t������`q>9��I$E��������>C�m��`��=d��,NJ�*��ͻ���g���C�\�+iJT���6T.Py�"f�/ ��޼�?��������HYU(*KS�V�\����o�W�����5��kT���'�x ق�dNe��xd��0��]��WFwe���	+I���#;�:�E���|�v6�_P��i|'�5�`i����Qn�Ѥ����=7���t9u���CGB���A�h��}C<�/�k�VM�]w8�"m�椣�!��7yVk�N��D�2	|=���rSJ�l����U��MT��s������s��})E%i��I��X׶Z{��T?��Q�O���B�%̖ǃW�i!�i��Cy{톹�s �����l��;�_^  ����y���o; .Fd#�©��،%�2u8)�߭�UV�i���A�=BH����xh�6�g���S؂���g���K�|F�C�J���Z�|X�����ׅ}6|�xWƍV�Cs�k�%�z�ц<�6f/�>��k(�=M0ց`Bs\�V�,�*�h1Z����sg�mCf}s�g"�W��4�4Ij@d(k��������
mo�^=�g���H����
����2e��h���jXnR=U4C��ǐ��x	������%]?ҙj#������4F���K2�哤�W�Ƿ����/k
W��<�\EN6�{|�I�/@K������]�����(53R1�/�I��ۼ �/�:���x/BCb���L��=�D�A<<�t���'פ*����M,�3� �B�5k����1,�K���w��f�(
vO�s�/��<�$��V�i���9 �M_Fʦ�q�=����ۤ[���i����^��&�A��xq�H�̛vRA��O�4����Ўb�G:���?����Lii�~&�R2��Νœ����G�H��M�3�����g����
��#*9+̍r�d4��-)���rC���9k�i�fxB1�h���Iy=��o�#�N;O焴��Vϰd��'Xk�c��~g �ו�pi3���̳�Vۦ��M��O?���k��m�l�~0<�*���V���uL�(�[Å\U�$�,H$T�hy�����T���Y�$����E�� <�nT�15����9y.H׳[Bt��H�xR�ϔ�f>~׊S�
�$v�bL�� j��1v����P8�EVb-8��V@q#��5^��W��o�o�4ns����[s4.�V.$�b�٢C�u���Pӄ�V�TX��.��J��k��e�hQ�J͵_�>���u�����Zꖣ�R1������ps.���9��Řo��(d�j��&0#�U�H�E��r�zƽ�ktG��U�`$�;w�:f��ӷ��=��a%�W�"��ĈȒ�[��
O���q���)�j�-��Ӳ��!%0W�ԥ�>�K�a�ݫ�%�����=��A�rO�X���
�[�0�q���w	>�	��ndP���W����*�۶a��EVR>����:I7�m�[��k�c~��.�M\��
.[l�k�<�p��,�G|s;F�:�DP^��DHf�Z��3ɢ�ڶ�_`�q2e4@��a��p&(d��Z�9����z��8�(��������ګ1�����0�D�E����#��yʞ�y~@�w���L"a�S���*A���"���ė3����Z���b���L�<�.F������i�FC�b�ބ7��~E_����@��<$w����VKˀ ��CB-�mYY�����~u1�1jT��B�û�
�!�8��:��V�����$SvU����=��-u!�)[�%q��r3�o����TR#_��R/�_Z�Z�ye^��'��U���t$#F!!QD6�k�=��y:�m�m��q��������Ҟ�� ��^�˨�H���� ۿ��M��([,t�*�Ξ�
�i�X�Z=�F�~1��aE��\�6��V��K\9Ú��X&�ve2oE r�2��,�Zs̘�pq����\�؊@5>�������5]`A���V��3�6�vb���e-9S�lməP���a�ֹ�ٽ���W�ʛ\��r�~���lةQyU�83�#%2Dg��Y������K�� l�� ��p�p� ���H��f�)+P��d�Ou'�Ї��D��)�X��B��wCU>j�=�X�Zv��x��X)Ar"kT����I9\s�B��j�eIwLu
c�}�s��}-o���u���֋ܺ�g>�[B�Y�˲P�Wv���y��!�NK30s��w���%�R�s�H���������ۊ=X!!_X��R1��~�'CŜEEP<dZdzk}���ӷ.��q�,����إ��BV����C�ցL�.Ơ/������sWDa`�9�$�DR�������\�3C㫔B�R�������/�%P
�.�J4k�������a(דTXkyUƣ(���%-oXO۫�)�$*��5R5�%��8f6�+�������'�0���,��0%t�@A����E/{A��A�m�G�\�(�\'�[ �8 MYK��W]�U;+����&Y�A��'/���h6��8�+:��&��HvC��{���:{�	j2d��]�Spy��0C��\�~�Z��c~�"���t������)m�˖z�P�V�j1����<�`8�#7R�~��B�r.k>�Nr��T1�0�9Rx�u��1�>�<���j ��<)��Ub�%�80o�3p����?e���T5�^�;����3J2ξ*~���X�HL�#3��9mC�K�����b��ݪ?���u��nc�~u��E�S,Gk�1^�;a.ɚ2au7Y�/ �Ю��d���e*���렶� ��OX\n#*�~�EB�(G�6>��n�	���L:+l�գ�'�㔥ۉ�>N6'�����X�K��I��Qᐻ?Փ%3�2���7���VU*��c3�6�NP�#����V�	|�{��o�4~QՐ��Q/��+ѿ?�\u�Tc�ޱ�y�h0E ��U$>	��+�ߨu��U���`/�"p�K[�[�ZAS?6��Ó�kR��7��4� �BG~�#E������n�j��:� ��Ћ�m7I7�w�֠���b�!Ԥ%���D<�	]rX�/͑�x���J_;�F��D0<�rC-���8���M�\�GΤ�@�-9�|�'R=6�}�����|�@U���,'�Z0I	�<�s8H4�����G@�̎ڛ��U���a��6����i�(���M���j�1��4��T3rS��?2�K�0U�G.m-_`��K����������S�dt��h�?;���X�N��d��&xNgNJ��^�$Oj�@��[���v�)3-�j6���T�՗w�>)�x��c �~�?L$j�:��X���H��m�W?~>Sf2�Z]�����F	4_N��<��Ku��f��U��[4���$e���h˰�'��B/�Rè�$s#g�;[�5�'poQf�W���"Y�)F�yU°��@l�;���1?�ƃc�Ħ��{���1�k/�lj'f%)�Kb(q��=w�w�<���.��\F�63k��܈�r堿bs�?�=��/ 5�0W{G�]���l��������e���cL�6�`�3e��y���lC�%� �ҠZ%��J�	���M�@�ރ�i�G��aF�vD�!���oQ���
��XYk��7�_����V��P�).�����@?-W�\��(��fW����؃�r�p*1ǉ�N�J�e�H-�xo�m�蚃���~BX�������X�����dtv�Un.ݡ$ު�1��p-"��P�$���wUou+�;��ʙ�Wr 5�(�����S�Š��zwb=bٶiu�a.u���;�^%��;:��N�e���&/n��'
z�yK)�o��/��k���I��v�R��\���ciHA&W��@|�D�8��h�};�]��
@��B�l�/qt?��ʧL������/��IJ/N׽�@5,Q�RVO9~Q(���H\7��Վ�*k�I��^��7:w�/e�d�w���%�*�|z��+�� qݲ��^ȑx��Q5����xB�S7I��V<�ٓß �dK��Wq82�*"|'(M���\��"1��O$�nj�]8`57$z��(]A!h����I-�q��M�A�r��µ��T�����o�MB�Ϻ�)n������1��dEQi������S^�oZ�x���� ��A_D�=�����{r��;7=���+�� ��BdZ������ ��O	�p:!��՜���������-�9'�Z1��n��o>�A|�֟�`��Tq#mGc�/�q�#\�&?�*s�ܽ�"Sχϡ�Z�)��+�#�(dΟ�rbjÁ�H��Y�� ��i�=�*�夗���){ʠMɛ�M�Y�g@4@ԏ�����l��oVA0�T4�.<��{�������Ͽ.��G̍�?�u��U{�ST���H>_t`.Y���@*Pc����s�;I�e�d���Q\H[�w��pǥ8���'5kb�k��k
��{U!�᱅Z*
��>��g*@034S�ӑ�Qf����Gܵ�=N�i�s(�A�0'~�e�T�[9���݆X����+�T��ǡzh��D�LۇTa�X�;Ͽk��r���7(�[vU��7X�2ʒ,Q��"�;��e�A�����c�	�C�1"�L���q���䟟0\�+�uZ:<��}���ߍ�Cۚ��$��^�|.r=BSWH��1�3������`���:��RY��_� �RkpϨ*�;�y�y�zt.��,�Y��n�_���-��^�c�T1�B'�n��◩���&���SPj�Q�2b�����	:T����]�s���.%�Y`m�I��}�x��J7˱�
q4#:1,n[���8'�
4�S�u���k��[(��{�ń�\����Ù���+�c
|��.�{�U^x�j-��������#-�7�y�C����P��x`���`�m�t �d��Ɲ�~�_O�]���$П�����ݗ! �"2b�~����4�"�#r�!��L�cbDk�:>��+X#�4i�^��d�x��t?�0�{�l7���\l���U����vޤ�=����g�	pU�������C59|Ѹ�V1�Hl�����鈀x�޺��*^  �+� ?�d�ݒˁ��3���LE���vŊn������n?�_hJ-fTg�~"+��=�vJM�D�eVT�(3�Y�&uKߤ�>'�q�`���46���wU-ҧ�/f{:J�0yЮ�2A}��p��Y۶m�Ϳ|�D��/}

C}GEv#��:��C%M%�����ۀm�8M�O�Q=���Cï��'�4��:��z�K�[RI�q���z㽫Z������V�yB��O&& �E�a�o���$��1RZ���O���ƅF\I"��sCMh%VT�*f��)�.��h�٬S�S�ߍ��/��%���V{��7��qȻ�5D��"�nF����?�����$?�窏~C����ԁF����F�4doj��C�J��M����?ĳ�S؈��m�$.��*��c`��w�*^Ŝ!��IT`��̜닷�.{�����|g��G�1�ѷ�Lv(�^=_�{&�?��eBX��M�Ë#����gv*����B�+�|i�H�j�T׼8�B'Sr����*6�OM��Y�,�h�7����'�w$��6`l�7�?�y,�i�&�������T-�&�ExX����]�S�ׁ��"2X-��I^r��a�ť�K���S�[�Sf�	��n���\1{���G0��I�(�S���-�F
b�C�Ў����xPOg{� �.�b�a�̓�P��܇n�z�a�Ř9FGv��P�sUĩ �{��E�@��ǟ$m��*S���.�,
��g��Z�澧Llg�0���U�> �X��Ǹ'����%�����*��q��_V����ϔU.ڜ���QTW|�������G%[f�8;.u	�M��_F|��Y���U��o9�L��,���ɽ��(��
�_�����P�2�p#��׺��j&ͺ��^��b`����K��}KC�\�Ӌ�ø�N<k�1z���C��B���"����+fX��x�(�[��zn�sh-�#J��|��p��+�F+'_cټ^b{F����<���X1�q�z��]E7�`�Zt�L��Q���
Њ1�����cfIr�c��/�_Vcޛ�y4�'�1��/�Q��1�����.�ykᒬ�1��osy݆���Ɛ�(~��5v�h�!K�'�p�C@E^K��j*�S��x5I��<�@��Q��j@{�p X�v$�pҧ�A�ݲxKEF�,|�Vc����+x�K�ߙ�G%9�g��*���@]�V��~,��-�/�f�[�-�� $+W0�|rDȨ�<x��y�@�_��T���i�d�����s۪���S%�#�=̷yY�>�a&�ҺX��X������*<[�we=2���^/a����'���a�f��Ft͒�ב#*�����t�-�j�g��W-W�-�=�m�WU�U�ɐ�Su۲=��<w	�U���i3��'wniѮa��(n��;���b�)8�A�7��f��B H��E��*����W�]*��¾��A��D���r�j�xg�ai\��f(�&�E���]�t� �����g�0:�&u-�9�+
�څ��X��7�&
/�*�h�L`��������h�؄)�<4�Y\v++�@w�Z��-z�x�k,�[A�)��O�L���\(A���c�b�H�%�k�S�PY��|�Gt�[Ajs����5��hS�CH�����f�j_v�d%�,��Mnԑ����+W��XI� C�� ���W�`�FFR�&t�t	���9��VJ�Z�:0��E�o�eJO��R��x.]�F-ޟji��A�\�����՜�g�%�G�:*J�1����N�`���F���a�)� ��Y�,�=�+Ș�}�j��*�8�|�9D]	LtٳQ��q��>�06f<����Bl���5ـ �:%(d�[����՗������g�{n�^��krs�P1����n�����A3�:p�RY�L������ ��tK+�wP��F���1v��5��k�+]�[��ws)`�Cfi�"� �u1u�[$>�p#�l߹/�U�T,�W�䬹;�����KR�����`�Wq�[v�pՑa@�¾�I��X$Q�УN����ˇ��`��_2|����F:6/�')����YC���IR� ���<��M�6�dGx�̣���h(2p������*V�-��Ŀvk��@�;��<	lbd�l�O-BU�6���5�b{K�3�{=|����DYB>!�\��t��z�ҎY��G�C5��=��Y�_$MG3���-�v[�
W�µ���[?�5�P	����V^��p	�=M�"����f^�=
/��d%��%�/tU��Gt�Kà�ȩ/����\�̹���ZJ�P�}W.|�)���~��_�}������ޮ
�6�i$���Y� ��e�����4y�Ҭ?�X���կQ>]^&�Ƌ�vjTŐ��	�]1FQ�he lM�e���4'+'U=��BE�"�����S�8���V���֝�gA��$q yG^s�����J��E�Կ����ۖݛ��yΩ�|�{1}+*�C�.n8��;�[��3Qm6��<-V�j��n���1l�i�H,��b �E�
�]��/��S�K��|�0�_ZW����r�'f�ϧ�3�i�LM��n��\C�	5��/eI�_Yl=�x�%���& a��꾢������F,f����(�����f<c���� �&���<���șY`��w��)�$�]�l��C�{��c��s�$�n'�������5�n��w��Wj�}r��hx����츝����0�l�|�|b߽������9А�6��5�®%��9.�
&��^ykhȿ�!A��bK�����3<uBj}��+��k�|*N:i�V��ў��XeEt��+�ص�	5#�.4;CA��}[�c0���{��{�@�<�t�:q�&�ɺM�� (�����^�s���g&�k瘖bv0�k}�ܒ;R�Ď�l/����	Ԓ�{"����`��|�
��	�B#�z/�ۄ�)�!L��WKow�P��6G�a���J�b����!(�#��@���G�fw�r�S��M��c�:vv�`z^��Zж��]�c�ZDX>j	�իl��1Wl.��NO3"*��!�3|3�}�uw:w�Г��\\)��i�h�������o�͝q���j@{��;2��~||VG�7:0s��C+(���Y�~r��s���%��w� 	�$Su�sg+�� �I�.�L,e�� �G�Sg��a�6UT-[��-�0|&~������E��o\C�2��<E���OA��ʭB��iM�=��avxa���w�[��>�H�-����-K�)wu&I��\��z��Du�����gs��?���@hl=�o�sHw�fz��z�`A��&��[� >��#F.jA��ܛ��t�m]��o�+dRV+�Sf��q^�̔r �6�w6.P@�t<�W��$��jm�ɒp[B��(������"��+��~Wpi�`�N���z\�P�A+Hj�w/�W�
\M\ ᷞ `ۼ�3��℺��e��}~�������R@�Go:�<���~O$�q�а�J�����u>��;0���} ����-��c
���.���3�ݝ�*�L_�Tdc���(v4��	��T�7���h��$��[D�ٝ��E��'i����C(N�΄��=��%��B��ߡi
LP�Q�F����	*-�*���yq�s!�F��K�^҄��s�}��E�
Ns�V�%��`���nf�]�^��4�����v��J�{`nբf>���a�Ŭ�a}��͆�5>M%g�ΐ��F�7�L~��7�g���T�?���c&��D#bEȩ�I�&�}����6���r<�0il�	-ci�Ȫ�2��f��r%�,W�L��\�oV�g���\�(r�%���	o�=���Gf�bz��������ڋ��$i��_��q:�t��R0
�#���t
jnC4�uآ	'^���YQ����2�B���q�@�X��T|�Q��~��"ΏY�Ay�TT��=�l�<�����Οq>���pc���ݩ�L�rP��_�z7oɪ����CL %ʌ�'�`�QH���z��@U�7ep_⧩Q�>=������ʩ�P���ޏ3�Y?����Q{E�s	�I�В���QCS6��#w����������w�QW|�b�tZ�/Iגۿ���?�$�^UuP�k�Whp��/�9(��VV��n�W��-��� �C�h�-���LC�����(�c�Q0�Ӭ���
ө�~��RP��t�ygk�͜�9��\��j�+�Dv��8ۙ�%�A�_n
�8�A�{O��5��� ��L���
��c=ˍǘ-yA)��P#%1uh��}W���O�Ip2(���g�1%�g�c�2�����{����nX����죋�����a;�v��q9��Tm����f;4E��G�J(�ړ��А��0�+?��*�w����h�]"�>DuS=;ʣ���U��}��E9�E$�r|3}�r �Ip_��'Z�@d���ꂮS5�{�&#	���7����|pf�F��C�R�|/
���+^�%)��K���X*�O���B�l�x�mJ�:�"d*}�t�]�W܂�:�
�w��� unOv1p��X�uE𛦳s�����.��_R�s�����;�jg�h��+B�{_�0�.�Q�q�>LPNs��ЁHS~_X��{z!y?MHx,�TE�~~�?��{������S��v������ ��)�pˠ�?^�2��㌛r�NMxV<K8��9`k�"���y���A]��.P"ɞ3�ټ
Yf�ü���}sa�.y���$��b$��pO#�Ɍ�1]�� �>A�DѢi&H���ܫ�\��nHI�Vu�vu����d���>0f��W`f�{�{�m�� �J�ˢ��i�@4^a8+�IA��A���b�B�tɗ���C/ZE,�yi��Bb��N��X0�V��Y,��.V?�R T��?<e�0]��	q��0�����H��A�Tc��2�k�͓V! �C�{����w-X�|]�S��{�P����σ�y��F��"��B�2n0�/��}p�^�{��r��^і�6}�6K A��,����-c��
�w�QQ����
m��
'��@o����x�bU�{�H�u�����$���F:�Y�gW����L杜��kK���'�
������T�k,���1D"o��Fv���v#^e"n����N��RM)��6���F���L�QΜ�P�J�]7
kVM��>2~�r#�J�����2J��P�V�ý��ǵy�0��D>Z�ѺE�jxC�3m,�/�ī�?V� 8c��� �5y�G"���{����\u520SJ���a�/Ƴ�D��?Z��g����� 8TBV7}m��!
y�A9���᣽8�J>|"��}�5u[��u�T�5Ee{�\�ʋ@d��Y��C���>C5���4�A���a�*'~���c��w�;}ma[�^Yv�����"ql��s�6q���9�KK�h�z�~� ���'��mֻ�:"�}�1^7�;� Q����i`Q	�g;�P�iІsw���zn�&����İDJ��'�����e^�'f�?��h�8��C;N�5 nTn햶4%@�x몓3gʃ��t8��*��(���z�u\�T����.vn���D�0!�3e�uΙ����qUT�ؑ����#N'�(ZGz睫� I6�#��e���;���Q�ïԹP��4X��P�L���{�v�b�\��8�0+gu���0�O���=f�]tZ�9l��w��k��To`QM΢��ؤpwm��b���
\�)f(̄G�k�m���;�z{J�����,���a:�Ņ����D�| �u�؛4�Y�5�$Lm9�CQ��o @O��f�y.I�6��R�T2��yuS'�Q�u.�D���]K,�Y*1Ua.U�W�I��e��d�}���mNZ�W����9,0��SM!�Guz�C|�QD�o�pC�����
�X�ї�%�G��ڕx �^}�3�(��F�y���loЫX�U[@=��S+BO_���+���bӭ@��$�<7�Ӭb4�z�������r�cY�'�T��<)�����ˇ@y���o�\�N5C�S�hj�;�CDl���4E��9�w��� e�=*3�>|��σ-����ur�өUQt)K�i�;N&�e�IQ��<�T�mU��G="���_��]T�z�޳8��m�?1��s��O��"�c�D��Xy�(����/+%�1�&�v�<��~E)%���`9�(�k���y��<�lR�;²C�CF]��W�F�sjD��ʕ��"[ˤյ $\ �@�Sf�E�B����Dn�����Nfm�L!�9��|k�L
r�ŦV��������φ7�����4r��.Qr��U�s�q.���l�a'����3"���`_lXz���2t���{$A��EX��'}���B�����!ν?c� e�!@jO���7�8���p��$�-B�3x�ND���pь����66��U��s���	��9b)�#5�P��2s_�Ѐ���ʎ/f0Ն=_���۵�:�+mej2O��d(:�!�l�H�dANoz�ž�"��x��=|n�w^�R~��Q��c�c���T6�3=v~�	Ъ��"�[?A��	�(}�ͺB���"�eq�yȅI�����t]���ކ1G�D��`imɸ���(u��@��X�ho���x�)t��y��f�**�{+6�������>U�ٟ���W_
c��-W*IΎfZ�(�7�S�����G&�j2v*��.��� NSꢿ��U�Ո[����X������n�Mbԫt&���+��ʖ9�t�}'��>k�*��V
�q`���� dr���a�u=����hY/��"�L�5�"ddK�y���ɖ����]�;?�B���2��Ա�h9����_��hFU�vZ�Gi���L�L�ᄰd�8vV]����r
_��_�^�XK�����8r	��r�=�,#��q,���Ř�G��s��ky���7׽���.��M0�?���䅗��jǽ��������8��F��wo��h�8���߳�4e��V��̶J~�1�b.���[a�0`1C��Bz0�0�P�xU%���7|z��e��"�^	�P/�9��	��b�ʓڸ��mS|e8�D�![o�n���Z����
",�l�'�����7ֻ������3�ذo��\70�?�DMʫ��Yx�DxZ��%*>����� � �*�j�p�M���%�B�wY���Z��f�bJFo�j	��e]�� �]��O�3��������]ڲ�?4�bpx;�1��`���&�K��
������HɄ)s9�?]�|�RG^5�ߢB~�Y������G���7?��b+Q)	ǼϺ���@
&3�>��ѯ����/�H�E���#p�l���{�'NT1r^��x8�2*��4$���r�&e���/��A�$~#��ϛe�y��{����  4�����eD��] Nr���+ ���X�Yi����%� ����H����j��Tm�L
��:e!�֮�rͯ�=%���ꡜ�!�X#�����[w��9jj��ˬ����"'�秌y� ��į(d�s0<�Ԩ}%[׆�!2�^�E��a�K��e�y���z���Z24��C˵8k�\$Z�Xw|��'�~�F�P�m�*���F~����X)��Ɗ�o�vk�K�8O��@c�k�c��g���I60��(���c��:������ ,& ��H�:q��(�d� �2��@4k������̩A��5�Fm�LX kX�ͫ�i$�L�����w�O���;��:�5�L.'�h�����}���͆C�E��]��F����܂ő݀�2SG.��$2_Û��9�^?b�˃U�z�U����#����"=��ް���fHt�-%��	����Ҁ�?���o ��x`�q:I=hr�lb��$�zΏ^\qO|�]'���*8�T��$v߇��}�'o�d���� �^9�o�v�췈O-m�[��Ȣ��]��x�$L\Go��m��a��n�|�&e������<L� À-��W�v�&�q�oC��V}&�h��.�z�W��ZV
qdf�n�h�זi��Z?��z�G��>w������O���r���hTG���i�*bI�]I�»u,ٺ&��t����������"W ��EP�L��b#	T��1\
��-os�����ye�x�:^8�ׅs�k���7�/��b{��@kc���gy;:�E��dc�?]��/�n���2��m!ޱ�p�� j�J6�r����`�"Y����I-�~M�BF���((!��<�<lcm}�xtU�n��4	jq�N��n�i�S��=.�v⨜Z����)~�`qJ4�� ���E��jbX��E剱��vݓ�
�J��������4��e����Fu��}�z1qFp�MR/�Jh���W��&������l.�ߘa8)�De��vȎ�xvAl^���)t�~aC�^�)���[���_8��[u���뱲%_���\�"P�Uo�Pe-������3���=&�6��yM5����C�?��hU:��̦�����+�v9���>��D�[?�߀��X���Dn���d���ҐST�Kv��Y�3_	p7;�lr���y�fDn��	*)�1nI���(�p������-�D_��y~��S�?�B��?0�e	s0N)��TBbr�b��v�Ս��I �j��Wt��Y���5Ѳ��K~�g٘����|��QB�T��M?�0o
�x/�o����䄩fQ���^��>vX�1#�½r��ɴ��֣��
���Y_��#��d�}��������2[wv2-���"�lbɧ�k뉜�j��\�2On�C��4��?9b�_�� �fL���#V��A�w%��#�} �5�&�_|H�R	���А1zBٹ�aaz>�d>%# +?G�	ڧ˓wk@������	*��4�~� �H�9�Js 38�[�>�|O��c3h���수�$���D�i<IFǲ&�İbF]����d��^��JiԹ;��hs���0�F�m!e-��#X��d���B�g����%gFv�U�l��RW��=Q�e�1�>��+�|�'ڮ>>K�]����;�9��)FݟKE�yZC��ݽ6�`��W;ü�x�����e:|�nw�.!}x�e�V�ӭ�*���=jTX-w|#�o�՜�F<�)H\���X+'{�h�{��EXӍ߮!.$A�1�p�>b�˲�'YAu�@4#��H5Co���.ȇ��Å��Jr�T��Y�$���&���_�H����iD[D�VpԞ�i������3rNkt���������}����i<fbOSD��ջYpXA�#\&i��L�ݴ���<���p��.ٚ^��J8 l �Q�=\W#�O�PCg~J	[R͂����ִ\�˚[�"W�O.঻?7p����i�D �6Z}���};g�K�c[�-Y��}q��'��G�dΑڡ��b�EU��a�H-e)���O\[�**/cN O,�F��%l����Щ�<d�Dڢ�0��õ?O��#�>�Lkm3(n`����[�e��W�w�祉�8#�.�Պ mK5>��T���� ���Jg��+{����]��r�����`���$��0w� g�yg
�ذ]��" �LD��sm�6U(�l��@�ȫ����r1�Wy��Ia��򻵰�� ζ��#��B��J��U� &0{���2����w�>��4�}:S��Y��tx�:"g��us�^bs`�A]�x��3p�Vm-�T��ҽ����Ƿ0�H:�4~�b�m�X@��(�wJt~�h�y��,M]��D���y�ꤿt�|��X;�e>�����>�Z�KV��bw:���vqmy��$
�k���_r ChfMvO$�( ���o2C$zm��̙.T�fqyl�G���=�]��	^&�V���}�7A�+t�G��k�jSz���$B`u�ݒ��K�K/K0�bg@��v�֡7��{,�bf3�vU�F��x��M�<I��U�^�nlhDy���|��/�ԯ	�>��B��wa��Y�ka�O���tw~�5���|>SovV#�H	�__���Ĺ4��Q 4��{���pC�U�K4�?mD�Q|�e�*�:�@�o,6M���W�ʱJ���T}>�LȞ�x{�T-�F�AxA��λ'ŀn�]����x�����q��+j%p��UN|W�9�!�H�څ�������>���G��Hy(�8�%h@�g� =���<#\���c�M��:b�!�W�.]�..��g�%g>����b�ݱ�-ޔ�Z�`�G
�޳���;,ډV>�v�7ˆ���X~g�0�q[���KDg5�
F���&�s۠�@�ք��æ�o���LC��]?9R�I�Kۂ3�ń4��P����5���>��hy^b�4���!i?��{W�%d�?j�!��@>�@�>ʃ6��Y�7���\_�h��tU��w$|��k���5I 5����<����m�5�C	 q3�V�i\��t�����4g���|�Ǔ�H�7,�
wCT��o�������g�$���2���T��^m�:������N&�?�t��$�Ы����Z�;�{�t���h"��OI���P!���V�I4�K�E����^x#�@���� ��O�`lA3�g��yyM���T�G�C(�7)���U�k�M0c�<�l�̗80݋'x��{[��1n��yߠ��g|>ů�]��"�1\w����RYB�����Z��-#YN�U2�ym�%bU+��,H $ �pN�2�x�/��y�7c}F'����iB��m���:R�������|�9�ߙbt>��]9Vz��k���dq�X1�V��$$ Af��1�
�̯�b�%�`����}(�{O_멦�n��~;}7{&Aڄo�X���l$r�C�H5Yᚵ�ď�"-5�L���[�8���b��x��i'S���Zs�xwR ��7���lwm@ΈX��}�3��K���t����]q� ҇�Vx��U���^nQ�^Rf%|��w�.��<��ǞĢ��r����?�{=�U"�8�Ym_GZe5|J�K2�: ��;cx�%��z)�}A�c��hg��[#�eŹ��=��s�#L��aR�I|
����<��69H�+"ѫ��!���yj�7;�1��U2���|V8x0R<q��oF��ϲu"_e*�
�|����l�`˭�;ӏ���Z��%�ޙV��6�?����u�} ~���h�T����f	�]�ü�c�ޠ��٢P,� ���e��b��=�o����-rX��\G�-��(㍺zp��@�Q���Vo8zsSD#a��[-�icP�x��.f~����E�<n���2N5N:��<=�oY��4�w��Xa��b���=�N�R�s9��D��_P�Su�3˲U�ar\:궱_e:-�XT=�qr��ڷ��ޚ�j�N�T�7�_�91��~���(8��ށ�:i��s�@�N����~�?-s�GSF~w"%n��Ξ�JW,ֿt>pLI���_��D�z��i��w�o���=��������%K���m ���/b���cU2�~-�L�6�NAR��p7q���[e���3$��I��eu�����ͳzh4Ct�6w`��#�@�+ј�ŀy��{�A���?����H��9Z&��k����2�l�\�rW$��疌ј͌nZ�`��_m���sw)�H�#��(3� ��i�s�(%2a}�W���(=�!�����R0��˨1����m$ݖ�r����v�����2x��f͛>|����R&'��L�.�����p�J��J����+��0���_��.�cQîs��W�i�C�qq�r�B�^M�('Cϋ��=��~5�&	�ГҒ��F���#�BP=bl�%��^��>]?Y˛Nw.f灎���F!j��G�n��8�q����ßH�'Q����~�"Τ?�p�����v��7�֢4ɑf\�4�X�r3`�6��զ���E.�=���?��N�!��T�����x��
�$;�ϵs�$���/ʘ-'�^
?j�X�F���Wr�C!-�̹�[�fKgU�]��9�F;����'���N�A�њ6��4P�Ro��ұ�ƾ�����q:V���B�A�d����!���J�~
��%&�y;v�X��*X1YO'�j) >B� ޥa�!�H��0���!ߨ��9ɞ2�_���;���҃�t�0f�TY�$Ƃ��]F�XN��.Z�|��ʤ�,���m��k��q_��)����ә۹\X+��:|����ش:{�H8)���IHIZk=n��K��3H˨�1:�<�uBh�1�8��-M���q�:����5	M��X�:@���U�Os����Y'2Ô86l���mE�������[.��_ 
F�?��zE"ei�.`�$}|z�:���JN�F���gw޶�*�j��\D��<gx�v��8:
Ϟ,Z(��j@��F}��\�XNA&{y�l��,����I��Ћ��hK*���6q3[��.�]��0� u�\'�1���LHy&���r�v���Ǖ���"cR�e��7�h��{#��N��j���$���MI���Q��j���W�¼/!�C
�:Y��9�3n�9�M��!<�z��A�rC^�#����/Y~q� p	D1��]�fo=xX`��i2<a�z!��>]�e����1��3���b�J ��z`����K�3�$�-}k�_A8���5�Z��l��a��*^��~�}k"A��� �<�_Pa�I 9$>O��?wW8H4�7Ш7:r��������6`;GC�X�>���h�&�4%����<j�Sij�tZ'�DR�O�yg�by�](d��l����3�y+�F�c@�dX���^�%�k�\e���˜]�����W8�ס���Q�7�F�3km�����?8�	�������]�������as��==)l�.F�Vuz�X��]�bj�QK����K�x\>��,�R.��+z�ϟ���_('S���yY����Q��N&H�T�pT+�sQ�G9[�Td��U�����,���əJw}X��w+׺�.v+��(8Q3�;����Q�KE(�P���l?֓�%�[Ou�1 )�$�{�͡/��߲���6mW�'b�oؖ~�9�?�<=G��Z��Ž=��a�.�Ll�m�R�Ԯ�=��c�-#���ۋ��������+i�$/+� 1������d�2�9ZX9[/�/&E�����c2A��e�L17q��$/���h��2}9'�+�AqD�g��Ԓ���!��g|nu��S4�K�~��k������dV�^W^�%f�7d�~�y�	����'�'T��#���͖�*s0i�:����s���V+c|<������'S�(p�=H�x��?x`A��&����������B���઎�z���wW��� �%��2!�P��k=�%@�����3�S�6C����H5se.J�v60���Tz���3���t�1t#�>���ڮ:�?����nK��ry>*t�U�j���r���\JY���S):U�N��O�:&{���s��������k����p-<Ӽ�;�Q2�������"jv�r���\�X�7��`Y�i��1��L�S���
�JaP�nm�'���[��ep��iw�EGr��ՔNX��	TQjf�o�ͺ�0���~�Pi��xY����#�GUˇ�]:�����&/+&C��vn�H���'^����4_�]&�l�u�MY>P��t'�@���ّS����%�xp
H�)�3���-}�HT��C��5�+��B�������×�@`{���j7b�`��5�8���W��{����6�F0��_��=E�)a
{e��wy�ĔgඓӋgg�Ձ�'�J����i�<
��Ҫ�A+�	�-� j�q�}�|��L���l����F�^pr�����N�	�bn1|mxS
�O�Ժ����Ւ�V�� ҟ����t�������Y yQ�rk�d�p�0��dA<g93$8�E�`�1uΑm<���rU�Ŀm���ݴ�L��l#���,��T�XlEF�!3�����~��w�\_J�l����jc�:�b�<-M�r��j�pH��_^����4I��B�e@(� ?;!@1��#Z�#ܪ�����K���e7�/�$�"*�wD˃�^��C�*:M2�;-����Pk�7��5	k�9�\/zr�4'5݊Q�'��C ݤfR���K��l`��bY
E��|�D9��걢��E���+� �Nc����>-��d,qq�{]�/xЫ8�ʰv0�Gq�Zv&/�/�	Y�$̾�z��T��	q�0x�Hf�s<�V��B����hw9Ncn�LK܍+�a|�r�_?Ɗ��o;�i�X��I��6��,��j�~t�G��{��a|é���]'��(�����E'08�6��OW��u��#�[��s�7�V��8�\��ST����lE��0�D)��B������I�⟋��Wxb�JQ�����Z�r��J����3$�L��Z���Z�"ޣ��!�c�c#��7"�OB��9�Y<��}��,Q�c[��诪z��������.�c�`���T���m}s�R���ďl�H�l+��=n��WܧH�nD��&A���˸�R��tW�l�a�sL �YW�G_��_�VmX�ۿ�đ�	�d5�U�c�;���شh�Z@���	��^C�iq�}��8�W���6�t����?�ы=�o�ԍ�`yO��*7�Aۛ��@dO\��j|���v��(���%�o+f CB!�#:�S%�Kog� �=�y�]@����p����AX$�.=�m��$���V��^>�,X4/������.ҐՕ
��A�3ו�Uy�?-��7���<��4�i���Kg!�O).3N�خ��s�,J���f�Lk��N�n�\��
� �0\&����vX��������}s��xrD���U��{��fLe(�5�@ܔO���)#�ޮs��I�;:�Ⅻ���\�f�jz���X����O6��l%%s*u�J�_T��5�Q���͎�A��]}��e'^�����y���Z��G�R�����&��	�U&�5�T�^M&� �����!�}����F���h�oVv���8O�ыՅ�+�zbI�p��*g3�9�a���������u����	�(��r��i�@H���4����K@�����^3��	wס^d앿r{�1�)}�?/0Q�.�)=R8��ܱc1Gx��a�~OvD���K�I+kJe���ڝ��9pxE�� h��1�fEQs��#f��ʎ	�SY����x��U���V�6GVj�k�'#g;�N����(����Ѻi�\�0x����F��7X���l�ԶF�E�A0�6G3K�͡5K�����wAT?6�	Xq^J��-�h:I�c
ǋ�xo��>j.jbG��%_��Kպ�ؘSQt~\���ݰ�Fo�aI�;
��������F�Z�,G-����ܘ�}������:.z�������)�C`����dV�S��;�92����������Ĵ�Zm�hŇ}Q=b�_Q��΄b��W븐h��k��6l}��D��j��������Q7���p���!�d
�8�zu'���|�n0pp���#E�zڨ���ٽEf�x�99&a_^O����vߜ�1����nk�����c��ZN"��tI2���D($
�5ư���C�z1�~��:%���z�o�	�:�e���"4*�y���ޟ��U��nv�DĄ��s���߾�����D�:��2��c>�<��i�	'zW�j\�W�s�Iq�\L�I�1��+�'��Cۉ�6+V���jʴ~v-����"��	�F��O����k�����F����/����b��1e�� �o0]Ë��WnO0v{�+��E98�3�̚h�؟��!���h���|�| �nE[����.v�g��=؁h���ɠ@�w���A��Dڨ���MD���FUg�e���k�ޡ��C�� ��P)�~�޽�І�q�)L��J���3j��1k� `���ς�z�
ϫT�,Cj�Ht'������>�\�����Cw6�~v�_����r��UX�z0X� �95˷�������^F*س�#Y	t0-.42{	VY�Jm�
�݃�]��+)���0��,vp��pXa�t�4�2S�W��%���Eě�!�y�u�يU�hE���Q�� I>�"4�B{km�ED��f���C�d�PY(K5	����WMR��'� =��\r\�`Yb��R=���i�	��G](�~*�>�a�QߞA�s1"��X�<l���*�@�������x��9�2�tY73�FԌ�:�4H+TC�b7��QG����@j�E����a���MaѪ�g���aAi��X,�٨���=堮�Bܷ�)��5��*40��V�;j�*��8��ĕ&*�x�w� ���E��
M���v��1��E�)?Y�C���RD$�H'�,�����ƭ�i˱�i�i�o �D�4pp��/�M��0Æ�s���f�[2kz�/t����c�p�&���?����x-���_�BA^�>;%.Qգ�����E�W�d�Eh*@���<r�5�"��0���Ѓg�������$�� ��D�esN�����C�r>	K��Wu���lp��3鷐~� t���͡Q�'Tv���Ȩ���^K�C��՘4:���ecǛ���.�H'�����๭�����SE25�,aH�]U�]��B��'�L?i2��pkf˶e�C"��|�s.|zXL��VI_`r�jg'�b�*���2ǚHۈ���edG^kqa;�Xu��C@��������߁�����\�O%�J�"���ji�8ca��>%[�2��S��{����`�JaW�F��$[.S "qΦ�Nc�Zʯ{�^#�)�Fr4�¤��*�#��Շ�}>�UZFT�@�ص��!��tp���^��UEU�8!J�ѤԄb�)�F�I5��y�h�'��+�8���>K���*]�(�]���eD��o��]ƀ����0� 0g��� i':�
���c�ʹJ��/@�{��L����`��M�J�;�7Y�'�ĉ��"���F��<�aQƏ�#Nۙ?`b��"@�"��]���f�m���&a4~�Q�cH��%����<��n���᪞F8�tv�x�.Ӄ�E�u�z�)r����m�6��i��i�gWs���TXN��+� >7��n�_pf.f�?�p�h����C����P���g b� (��%�������QI_�{�2�v���t�gk��I�!��)>-z���'1�At��j8dys���!֙|�qŀ�t���u	CK�	��^�M��!�1��a �X�U>��B�`�Ax�V]�.w/�޾���V4m�Q l`����ر1�(n������m���"a�~�[9P4���S�����+��@!���8�	�&)���t���pY�7e�y���.(B-�^%���2��N\ʹ~6�� ��񰁷1����6�7J�M�� 
�̖-�-`�rN��7Q��L=Х@��\R&��i�V���������ʉ߷X�-�E�~�=	|�o)�w+�S_�C�}��W,O�Vs�7ΕS�F�6�/�Њ���;l#��b��HiY�Df���j	�΅蠲<>��c���Q�)�}O��7j��_WB�	���x*����zЬn�k�C��"w��)���(��U$���
Q��[8K�|_��&X=Î,�i�8Xǭ9�������)��f�+��>-8�L�3o��e�/�����8�y+�nԇ3�|��_���g�̪S����%��U�FS �N���N�k� {���g��;��$W��ў �F,���AGl�	m����)=}���d9yc���t���+�uRx(�	���s�姒�n�7�9+���V�q�/?�F�W�V{���)I�xr��ãFƲ���3b������v�"��r�q��*��Kٿ?� C�2���cj��������^v�<��py�+�^��P�����u&�Zȉe�UP�T3OV�J(Mm�����0(�gO������J��SH�d"wcW͛�Z���$���҄��7�D��+�뺞h�M��En��b���ǽˡ�`�;�D���E:�l�A/)��_�o�j�$d\m��d�!������u�?]��i�eWh���Q	�v	M����o[�s���;vm}{��+��[#�E���ȩX�����W��J�@U�?B ��b����a�^Cr�|�@&=��mj$�>X?xZ���dXx��A���=$}�ه�=�0;�NwW+��'~eU��4��4�/���G��h� WC� ���.�o�ă�&�C���vS-ڠ�8}� K5`��cC)��4���+C�JǜϘo.���ɚ��ȷ��*9y�pp�ky�Xd���Җ�רdS�v��2n��^�!��|��y`��s��F�G �7c����?��k�uUX��s�+��B�����am���w`��p{�L���!��P�\޲ޟ������XũQo����Xy�[U�@�r'L��L� ��<��>������b$��PC�Q�����qd�n\�C��.���m��������M`YG�7*�=/��)7O���e�%���A��;��M��c�9���7���BR1�Ԥ��2�c��	�ՄH�����ʞ�(X��#`-���A���1KI
�Ά�����ahH��(��3�	�
g��!%���
&��,D-����*m�<<�����TZ�x�����NΠ�?��`gw����X�哷�����ϲS��z�R�w6�ץ�w�����u�Z4�&�on�#\�� �E�����>Ҍ�!bO �K+�����ʫ^NPh�y�Nې�Gp����8��3�٧观BKه_+/pGI�Ǚ?���̹���xCډ�]L���\Q���%x���H��Õ/�2��V���4a��;,�geO���_���ph(�?y�I��=�oU���kR�QW�Wܩ�}��#n�5ڏC5����j����-4���ii�uYnc3n�����,����_�H �����	ݸ��R��\�%�.�y�d.oa��r�3�����y�J��x��e�v�8g��)�@����%Dl{�Q���/�rU���~&[HGgc�.��x�-�9l0����������Β=���EٗRs���S���v�طotȊ������3�5���I���n�����ժ[]7ѥ��c�q�Nh���A��S��L�+����+a	Ϲ�.�s�Yh6}��j��i�!B�\��vd]7U�ש�l.3|�E�#h��ܽ��q��#B��Q��'IWkE����q����N@�+�E�fl\�"P�-G�&L}�;�w���/�~���%yO�C�Z��#���e�H��N���|�w댔��sJr����+xZ���\��m�Vn!W�({��Zl�Yp�2͈%Fƚ��6����1/�b����[a�G��F<�=��{��y�C�Ɵ,h�؞cL,�|���K��j��2ѯ��<0A�ݫ��oU6:��5�W�a�N}z�Z�a��Ű�`��U�z0��?9%ev"AZ�)wh�&%;��,�F��Ú��5e�j������֪xp��m��9]��Ic�����1����L�<Ɇ��q�|6��9t����F���,D /��8p����j�r{V���i� ����-f&{#�e5p#,� �`GIz(@}��|Ɓsl��,l �c^?���^K��M��	�@vL�v 0���J㫔�>�J�1cE����$�b90���ߣ0��I�@��OL�D��G���˰��"�h�_1/3�!�D
�s��'���D��iY�S;���>R�0Ra����D}��C��y����a2Sd�s��:d�y�Y��]W�zU�Lf[���L4����*���'k���m����\~٠�����+H,%-O!���y"�ǖE��a��ݛcyxC4�u�*8p7E։��4����gѱ-0��[x.�)����`��K��,ۿx�ނ4���-�9k�jw���c�+I�ӿs-�R�|��+�p�������T��g⵵� Vm+��e��;0�o�W%�P�$�����u�Z�#G���ٻ;�� �
���5�8'ڱ�,#��8���QH^�7F^)�٦}&ޡ�4�� n��J>c�i���W t����8ٌb^�v�N�JK�r@9OŇL�.���4�Ҕ�{��`�>�אY5�4�C����Bq��hs����Ō���|7�hE䨮,��0��d�Yo��ӟ����<�<F�{b��� �"l��D�^�N��6����fI��-���p�c��C�XY�����Z׈]�ڝB�=QQ��&�Z�1��XȻn.��nKˠX���)n8����`yfm��;)�Q��g��q��`�	�cn#R-�X��.��s��)H!Wϊy�����cz.��'���g��H�#j��3YJ1c�C����m���c�������С.����&�i���)�f���h��Gp�p7�*6��	/gSs��x��o�u�&�-j�l{����0�D2�� �_`�\��$=y�H�MZ��H`���d�'�W	���B����#ֶ��	-�e�P�~DL<��nK���"�p4Eq*8�܇��@xV1��Y������lĄN��";��	���|���Rq�A.�-�TF��M/j;3G�w��ap��3�^6�"��Ɍ:��0�<ΰi����a9�m����U�w@��d��B�����Kc�X�[9�#Mˏ�f�> t^3�zI�q!�J���L�eDO�l
�9ˡ�vȺ�F�V���=5nW�-��a(����Ⅻ���E��y����rI���Y��Qb�~�����V�0������|4ݗz�Q���=
��2���{��x�%7x�Ä�Ź�1	��gĆ���D��������O��Xr{�f3I1����t(F�j,7q��n�KV�]�	�ix�]͞�4p���d���/y��nM�$�p�&3�V������Q���T�2q5�bx�=P% T����W`f�=�v�Q����.у����u�p�L�6$|VE�CW-�4��x�R�5�~���i|�[/Vr�(s�)�C���kF�*8��YU2Fe��|��6�#��.|&�~��9�F��
���&�l 4�J>w��U�1X9=��@���)�9j�"/|"��e
<7�˼��j^���%	�����:`6=�G*�c1����)�:[ P�`i�݅���	NLT��mJ[��B����j�xTR
�I�=?���@�7����A�a�}gû9�A�~#_7
�ͧX���s��c��-s����q��M�+�6��9LZ���F��^_���!�W]��%x�[�Ov�C�@ r��:�޾j��æB�4���s�V��-W8o'U�� �4]�)z�����v�sT%�t�?�:��gP�"PE�D=��b��V�.��?�:�oCMR�ЩU�fLa�������H��;�	�cl� P��͂���	�k��(44�c����6���8��f���ۥud4!L��u�+��c�Oޖu���?��q�ƞ����K��0�c��Z<�r[��Z�Uw��g�0�޵u�-��Ӧ��0���V�y� �T@S��`_������=��C�My���J�HnCŅG�'#����.�H�k�h%/�% �Uq.�E��<d4라+g���,��_�V�z��㷴n,h#c�''�v��_�lWj7�a�d��G�n��f���@yٌP1+DǢ�P0s쑄�p+r�ce:��RLé��T0� dg�D��������>S`����x�����]��)ꏨ��"�+e44��m�*:��+��^�ln(�	M���e+��s\�:�:g/�{
�*>����Ӌ�w��ƮS�0 ��  ���peP����Ur�i��%��<	`���O��+_rue��@�����Z]z	�Ulz��q����r:W�2�⚴.r>�� v��8��!����O}��%��+��9�
�o�EZr�1�q,��]?y[�?�SO\8�" 6�8h#Q�-����!ଳ��*�Zh��)W���%�z�ғ������È4���,���@k�C; ��ſK#1�-(�|y����CF>N��5Z��z���2|���^�$m��z�t�C��'��XKUE�2Wm�����@8u�F��q��M����0k9"� P�y���_I���T�9QQ񕻄H?+���Rw'js�~�^�gru�S$�<�9A�V�:�{�+�w��3*�Gn�aw2��9{%�k�p�o�d��Q�|�	YЎ���=z��x�C��̥�"���`M�3v�>��߹�L�"����:!��h�R䐖p̣�[��a��=fEh�5�� 6$k/qh��X�F���i� B	z�tgd�KVĦ��R{��&*�X|@�Cz�JJ��]|ڡ�%]�K��� NE.EuG�'��̈KN�P蚑ٹ�Q|��qL ��j6�-��3��Sh[��;�aз�������kB�S��\,���O�q6��jK�M%g��W"���سe[-C�թ"�Y�։hAi{,��27M�����A��8����贒UW\�Q4���2>�DgD初��=`�[q���S�Ɲ`���_{�D5���K�q�Y�@h�P�ж��'Ó�J��U%��#�$w���4L�!t��Ր}K�۲����Q��0}�6ښւ�&��,����@�V�5�)�R�(H�����Quc��{��ܤ\�1		~A�����6
�$����L����,˼2�4���%�E�$ȫ����r1ы����4!���q�����a@�8_a�
�VJ�{&��Ҕ�� tԾ�X� �Mq�n/t����.�|�0PJn	cU��Bv(�y*��x�������<��	�]����'�E�^������\�j�Jow����9g�ߍ�($���<6c<�|L���e���֨��V�gO����5�a�6�S��?_8(���Z��2��K�k����zOо�?��I���)������q���j�������ν�JŶ�1XH��9�쐀�[��][N#��ߴ��m�k���ܾ�S*j����5B������+����^�%Xz"P�����+_�P(< @�WE� J`p��ho!�k�u	+$S<�LEKΌ���RtՔy�'p��䯳�@�f;�`
%��N�4��+ߩB�A�v��CU"�4�3Ȉ�Zhv���84�W�3����ESJ?�7qG
�=���$��	��M'��s�;�Z��壔Ur�+����#�/3�%\�S�f���ҳ�c��e����n>�wo�U�:8�c^�y�'n�ܷ�d��=k����H����Z,����s��n��,��#�D���AB0#!*a�HcB�yCe_�3b^ΰ�:�A*��&���A�z�b`]nƚ&q�x�U���i�帘|�DPp������в��:`��;�d6���΍���ʀ�
֐2��jH�wx�&�O�s'�~�+۪s�}Y�[�0b�"�S!Q����?5��S�o��h�-;��Dd�!��CƖ�� Վ=���e4	$b=���Ց�!?��<��[�Ֆ�[�׃�28����M����_S��N0˾x�.���'��.�=��S&�����W�m�����Ȟ7	7g���X[�",�����&��y��(p���9�-�'<��m�v�8�uyW�N��ؽ|"��%)%`(�h�@&�7s��o1���[F�|U-;�xr��
����Vx��Ş���t���/kJCC^�Q�/>�H0�&y��w3�J�9����Y��;`'��zX�����Ҽ-��ƍ竄dp�]t;^Ѫw����=d�o&�0t�ft<��~��ov�&���{����o��X��imf��<\m���p����c�p�d<����LѩA�E�F}B��=��$5�uo�=�g�ȥ0�$d�pQ�T��Zs7P�W4Hc���sp�V�Fd~�7-Z����D�������e���&ѶlA�W�&LR1e��
œ��������\;L�=�%d�w�w����R^�4�l��v�z����û F������c�&d�J�:�s�&�F�@qL�)b���CjTZ��o@�{���,�6Uwŏh��$������A����ge�H�r�d7�F���ib�S�K�[,9T�
��(���ƞu�'�hU���(�4��8� 䍝�.��E�����Eֶ�Q��}���'})��$��aaCRZ}{����*9�T�k��	��(u�z7��.� ^����
ۄ��z�>�Ҝ@��X�X����|��{��j6e�� ��-,(X<��nr=��E*1��>t鑘���&����n��R������MP��.&R����k��^Z�p5�,��1S_l�B�g{�%�([���_ Ɋb/#}R���=�Fʤ�V�o_��ގؑ���$�Pnr����9��o)� �ÇLvRʠ�Cp�����&���\*�-� +]�T�R"�=�L���z�e�s����7bRC
�������!ӡ-<й�C֤��5��J�?ta:Қ,�I�v�K��50�m��m�ؒ�w_3>"l7��S�Օ��j1���j�Zbx�&�����q=9���H��]e]E<���荆��,
ཱུ�RW��	�K����6��uHo[�7'\r@�����8�E��&�FZ��˦�80���>$,�x>V�1\ix�иX��R��e3~N��?�lj�C��a�:��@U�B,2h֫��ƀ��i��j�(���J��%c��Z�`.r=��@u}��IΟ�
0�$�fYll1&쌭�MZ!�x�Ӏ�/C錛�6�e��=\��J�ΙDꤧ���?�y�J�|��������e��x9�����_U�����6W�^�{j
P=0�l�C-��8�Z$��u+�}�l��AQ7��t��gmAV�5���~��S+wi��XRP5��CT dk����u��3�e�r^�'K�V�m�B� �a��  y�!�Vez,|��TR(o�stN����3l�؊{�r�VR2��L����]�����"� K��Nג�X\0�]��O\H�}2��W�q|�<Y�a=��U�]� �R�����O0`���-�푄���r��#c|2�7�&���U1���7�d�/e�Z0��������>�{f��Sｮg=�9�ɹՐ�ў_�b����'���Q0LW���� IF���v@;zZ��5����x����@xQ����Щ2�`R �"����Z���*�.�JT
����Y�"���W��FD_8K���'F�G�|3r#����$1���#�	��	�8"'�D(=]���7����=5xgh�D{�)�� q��.���#���=k���c��N8� 4�"Yʅ�������x^�E�#	=��	~-��De���X[�M���n����c�1��{��$a�-�> �Ag���۳��F��ǫ. �_W^����o�g�Ǚ�9�|"��f!]�)��a_c���ZG8W�Uy� \q�pW��[���[�!��HW�� �����O a��B�x���s)���j���2H���ޭ�;o2]� ;��{�.�-U�S�T�������_ݕ8���O��M�ď��O��tL����xt��qT��M\D�(x�|��32��'	V9���l;�-���ݰ����*
D���&�2���He+���T?�@~Q�Y����	5�^eAK�?�;f���x���ŬT8�W�l74"te8.�W�t�|7�i��{�G����+�޷	�:\()����Rt+X�t�y�ޔv�!���
���T��9�C�9�8����A���5���:$3NAK�����)����j����6!��4p���]iԇ.���h�"�Qy.��W����7�����E��A3.��ֽ���g:ʭ0�����솢wy7���)��>I$�К �3 ��(v5q�2�TU��� ~
&���������n\���۝�����u�ڃ�������+�밡 �h�V�˟�þ1v��9�͚^����y����a�;��U����2�y�����^�w�����p�"����Àh>@7:�½~�.�~\��y����g�E���ȫ,E��l]qr�I�qEˌ�ӗe�Y���4��ws��"L#��A���T�36��S�o�1��>�]i�g�����@���X���y�j-P*C������羫^"�eb����(�a8��Oa���0y)��<-���ɪ���_�����3C�Z�L�:�ߘ���?�;Ԉ�����(E�8G�ם��JwGD7�|sX�d9�	����$�F�env�ξ��K\d.�C���i)���rM2��2al�ʚ�lF���z�?y�#��h���ðc��"�o� ��� �|�pQ�is�L+N�
+�e�C��u�:����:(2�����a8,�ܩ{>����w쓍ai�8�B��6n�  �����-��ka���vFjt ���r:<*�A��v|i:���8�u;��3���޵�������T���G��#��6a�Ss�՜�7�H�!�b F���>���H0,����!���g���u�U��S2��ar�}�c"9@Vk��,%WID}
�$\{���F��̀��Z
�L��8M�e	�<Ĩ E�3;��mG����U6x���)kk����x{A�j������O������4=P&�PP��"TW���BZ��]y+g2�/L�ӈ[N�m��Mn����]ԥ']D�Y%�_[��[�o� 9��3ü����ݻ����z�5e)!��Ż8��^��r�~���X�5�w���CK8�߿ig�ߪ�G3���.���#�Sϒ؍�7u�#0�����h,�D��X����X r�j���5S�H	�T�|�G��o��R�i�z�I9��{)���&3pObu�v%� �]&߾�ђ��
>��ڡ�QOJR*�c�+�<�d:"X�E���0�^/���Y�����ث��9��.A2D�������l�5�^2^Ԁ7-7Kv�E]�)���E�p{]m3.�5'^�G�~c�4�g��Ab��Jeruj���%Ԝ`�,��v����q����(gԐ؝f������/�&YԽV�ж7�)��:^}�ہ�@���l����<�`�������}�)���}�"[��}<�^-�^����pmٕ�ƌT�ˈ�!�dn��Fz���ʚ�5(�)� �'�)<ӹ�F3P\��Zیv�Y��r����T&#7J���0��2'�f�IzW�6螡�G���*�X�j^h�sT�JE5�D'����ޡ�Y\	Jrܹ͎����J��Ǣc'Rj#�)�g0����ȩ2�ۙow���WPD�N���y����a/$�<�Y��e�vrk�1]3�o��ZX�����`�7�}f/t�H�D�ٖ��T�,|+I��&|����M���;�S�]ˉ����(b��xkϞt��_��������*�2 |� [�_�l�A�����\�]i�ŖDFX33;5�B� �t�>���H��\y�$�lwWKF��� ��@�-��Yy�A��b��jz-�Fr�	��}v�#������6֦o� u�\�b�:B�9*8�|ӻ��?W~��)ѹ���+�*n �r0oQ����@�;�Ʉ�wƦ������C��GXg�#�+"���y�7b�Arr�c/������l5��T��P�R���l�����ڧoc�J��h��9������wKOxf\'0�v"1�B�GNK�D�VK�'����.��"��#�̛�4�����U��OR��桳�m�J�䐺_7�TE�c��ͪ�^�:�����:��3
�5@�}
"K��U�B�5ܳ�!T�2��i���b�U/1�~��-�>��iUN�q�~�[ju9�_�j˵���1�����@��^���(�Z�4g왪�E;��o|�k�#������gK��E�5>�Ӗʹ�?�q3��d|�z��0|[��$��0?K)p����wp�����Zv�{Y�q}���.�ׯ��n5��ź��<�D�Jc`P�v��zM���P��yKi㊘��e��w��%���!���z�����W6aLh���$>���/��*���^^"�J��*���P="���Q�[E�F�`b3��
�$YB���Ԓ@�A�?�R����rɰ���W5��yR��0c.���Ȅ֋d'}BN����0q��ߴ�"eS��п��!���8�����h:�q	l�l˲����E��'�k�?r���?(�X�vO���I�;3W�^�
F��0,j�Ϟ[pw� EA�&�?�-��Y�Ͻ<{S�G5��^�!�t�L#��'���
1a�S0��}Q(�,�S��
/��˸�a�V�`��8J~Т�T�e��������/=�m�\Ԙ��=��J2"�GR*��t�Z\�����D�ɲ�,Yoq�6u��I�M�\��>3�̩J��7���o_�WT�(�H.�Om�8�Sţ��������!�&��j�o��G�͚?`��񀙿�������
���P�uHl��[�;�=x�\w�sI�A���9L3䵛*Bh�?XX�N�i�A�2	@�e�G,T|iG����;��vEzs=����C[�./f�b�A����80\��}#d̑���	Q�@T��S#"~y�V��	��y��Ƚ��6�f[<��*GD�H0�`D} �o�Q�cW��g�	n��qS��ֵ�|@A���&le������?q�Sj�#�ڿ�*.��t�d37�"�]��	�vq�ψ��`���#�T=�Q�,v��[�v��_��@��b��=#�b��E�nUH/������,�׍N(F���N����t�!A=�ڃ,a_���x�+[n��!,Sϙ��Y�H"OCu�tۓ�_Bd�1���E�W'����ץ���:;w^�]3���lǈt��L�P��Ǳ+?q��k`�c��e�蛁��1<}�U��(��R	��E������a$KB���5��\B�[}ZnQE&�V��ڗ	|�c1K3���z�D%�1C��g���
�uD8�%���/h�oA�j{m̖�����
\�o$��e�a�;�8펋J)U�<B��>#�?��`�8р�e����=M>a��x L�K�pb�E{X��R�Z����1X�$b�˴/f�a��<6��)C�'�3X)�A�<�iI>�1�+j&�g�>�'޵'T��/禟vpQ	����6k�S^�z�����3ΩL�0�y�g[j<e�h�V��E�Q��<<>]5�Oj��Y��!I���̄4�No��:W2�]�Y\�3Y���9�(nAIP�͐NV}7�a6�l��v�Z�h��Q%��R3X�� �Rٟ\�C�vK��s�:~�R�xg���Ot]��@G���7�4_��W0W�F�O͂���?��w��B��r$R-��Va+*�Z%�%q�|�Q[*�/�����_º���1R\�M^`�MLW�"-�T����.<�d�S�v��a`V6����M����;�z����w	���� ���W���z��hz;="�W�X%t��K������?�JϺ<�V}"ɿ��G��4O�{�|�Y�=��I����.%%E$	�7��Exf�T�?���]m��]����*�~&x��N�y�|��T�#�4ܻ4��>�(\�ƨ{�z�1�������fĵ��<sj�oU�z8���MjR~�;��z���QI�ώ���c7j)������g�Q���To,�y���9+�.�%effᖏL|jh���.ݎt�wq8c���I�]��Y���T�!���la�C, d�f���&I��[������F	��c׹�k���}V�4�
�-z�e^:�`J����& ,��I���f_�����v�(k�P��"��}@XO�cr��{����	زSd�$ =�\~p��6>������r:�Y$;g��sJ�T_�<�ȶ���쩴�^Sj�'D.�`I�(  ´mk)Q�.��.Iz]^����R�|@��C�-p&�_�9�1<1&!u4y��ƾ�x��z�+��d�Wr�VM��%/�Э�:�y�)��=�q|VX`�Xc��w,Ġ�W�j�~�ֹ%��Yf����Mʂ��wrktM�}�Md�Z�p�&3`,�w�.P�U����CQiwZ����٤_�r��ŉ���V���/�j��[��B�ل�\�|���S.{|��O�$���oWC��6���������u�
R�����WDǺ���/�"Z5Ь7��$�1�����W��[�?G)�(�/ӆ�I��j�������̱Z9Mw���	�ae"��D|^��9ظ�K�Ci-��'���ڭ9���!C�Z�v5$Z�@�Ί���p���qǕ.�(7a ��ve�i¬�,��:Jf'��t����1�+ی�[_��s���=�yjFcoq�Uf^<5��	�嘽�6U��\OU߃��}N�	�Y��>�8����[��W>��.WV��@$�Fs&��|�7t�fy��T�����f#
1�H�gN��ײ�6��B���h�׃�?c�M���mn��?��Ѻ��H�`��8��6n�� �2�5�kf��`��Z���FE����[3P��H�A�0��)8�9a����\!�-|��
�wN���$�it
��0UɘkD�U���Ƹ�Y���T$2�;�`!VM�=6Q�"����$���ӎH7�k���/�H[%z��H�4�5S7Ȇ�h�����D�������E����33�G��gL-���[CS�DVu'���}�*e�[���S��P���T��1b��B���pm6UI�r�3��?�wJ��wSi��;�X�5���d>qU?3�����0�jT�u��-�]g-q�&�뾃���!�`x�Fv�ˍ3\�9���x.	��.+M�?���S�6p&r���n�,�w�8�`@� �?�_���x�`J$M&	�����RS��0����J��>/\[�3*�	�uБ�X�[�ߔ�R�U�[9z�R5r�s+��Z4g�=�*ױC�^a%�G��� %ae�,b�ҫ��\�azb[�����akb����nPF	RL��v�V�N����3�zCoi��ߖ˰���������P̘^�=>����l]n� W��s���<2�/�k�����G/�S��+����{W�C��6'qz�_h�U`@Q�#n�8W8������v-\�L#�|��8Jƈ��Q��%���v����p��?"��]���@�	�|�G���BX�n��B'ӫ���-��7�iC��y�%���&��w��j�n患!oI���Q�Ԉ�ZY����xJ���V,n�y!p]�=��f�/�K�y�'έ����7'}���h��pp���ܮ��v8;�ULw
��Q�vt�D�j�@�L�GH1�6HK���XUB-�ST���n�D��������-�t"�>0^���L�m���G�	x<��7쒽�)Wp�1�*�j�mNi	?�ވvq��)�1a� d�5q�E��6���SL�0VGFo�d��}v�Ii��Gq���K��Wd1$f���7F��I�9q[�]���;ލ��1y�׉.�~��q�`iMX(�v���8X��T���-�:��
�'t�����Q� S�^�w�.#R?��6�8 4��/,?lT�˔����q�� z�������߁�ץ��Lz�0�$��Ee�5����Ku���b|��`�q4���w��vzL4�q6(�kx�a;��(0D�¼���"e�9��0hv(�ͭ��6!赵��M�W��D�@#_K]+;��~K��y��	��c�Q�ѽ^b���`b��̃�����B��g�E���K<=�N����x���3�������ˆ�݃c�R��:����o�#��(����͝�ݑ�e餿��e���b��<a�-"?��@���?�|���n�����2:�Q�3��!�أ���H�ˣ'J�ɚ�H^����ga�_��J"�I��ʴR�t20_����g���>Z�l�Q�!��8ZY3������^�/�5�-�̤Ov�Ol�E�eO�Gc�#���4�%o�L�*���~��m��	��.��op�j1P<D�R�1	P�"���w>��$Rl����U9�џ�kDf?���9@��taf�N?�����"~�&����	u�u�j$��$(C�����f�4U�jZ����ȧ|�0�<�0>(��.h�j�a�KFP�����J5,"'Ɉ�b����Uā��z0�R���t�n�a�>�d~_L����=�Z�sr��4X��әV��=!|r��?w`O+�'���r|mءm��Ny<1P�T��5�&�#?+��������}F�G�tjtơ�oK�K��
S�}˭�F�B�
�@d������*���T϶���J���E�/ׄ��O|Z/;�fw�B�w��ALJj��qB�+�2�]��۫�q�>Tȹ�d�}p��!B����P�"�Ÿ|����e�b&f�w�#A��ZX�9wj�0�Os�p"�����ȴ�=C�o�?B�ѯ������?�|8>FW1��_.f�uN"r�^?<[�A�k�WzV��g���A� `6�#� }vp7����hn�R-;o&Nq{�L�U�%cr-��z�U mP|��DX&Ȝ��#���ާ�'uT1�Q���ڗ�C9jD�g�A9�mx���s����~���-����q�"���.�R�l�_7tf突 S��O�Ѩ���,g��<��3H��$ʚ2�.9��xy��X[����l,�1D�ޗ�[��l�5��M.4������^���{)��2(Rn9ڑ�-��SUÖ f�ϩ�<�~v�g�]�6(?A����$��-l�C��%�9c1|�L�[��z���\^�P�ÉʀH,9��U9��`s����VSK6@�����)hT�M�Ba�k�@�<�
�h������@��1�6���OZ�6���=&$ƢP=?�Yf�����)$�kaA����a�U~]Ohy
���V#���jyY�}�Y"}���j�՚��bn��> �"���b[8.�!��Z�0) �zXJ�����m�@���ۘ��]!�*Ad�!����i{&S���/[���z�W�$��^3�~m}���P�d1�˲kBG�aʬ�MHL����Bf��(�y�h�?.�Q��#v�ݰ]���������#ʘ��m��k}JW��t��;���M�nq ��Ǭ^�R#�DV{��[_ʚ�ކR?��̮W�0_v�!�r#iᶑ<��u�-ۢ,M�L=�S	h���>I}^@㥠+�~�ZRf��9� �{"+	����бxC7��C�é��v�%V�8����8��Uǣ\PF�����x�L�e���abS?�ME���[��1��MD�޲I��B@�����b7HT@q;�Iɕ����Йoƞ[�&���U���� ���ݪ��*�o��}l�dM�V���$�b��QL�IM��6�F�9&�Ɵn����C�Po3�ᮧ��Zw��P'�*%�nu�p��=���ƭ�WF��󟃽��Ց|2U���S�P�#�5�PAop�W_�؂�'i,"ca���Z�b止#Sͷ!�n1mƻT|D�g�A��oh�8�Į��f�~ :bK�ⳍQǤ�mk���֠�KB"�p+�f����:2JbkGK����<!�
c������'f�̘]_���Rdl5V)��ߺyo��#�R8q|�TNFݚ3ȿ���ͱ���E�>(�-�b��zz4���NX��H�����Z�M�w�P4Ҋ���$����zq�r[�y9U��΂�*뢱�4�:�2:�u$�o:��B~|�ѣ2i�xmV]��E��c�QݎBC��
��
Ǥc&��ھ˂!ȋ
*>��ɜG���N���䝲 tv�c1J;�H��( �;U{����E���<����0sܙ�Dn\o��Bul�N�b��#n�I�-W"!g���~!�C[���(���"�>�1�iRm0��cɫ�W����]d�ɷj�Ws���1n����ۮ�M$��ّ0���j-u�ּLV��@��r �F!{)��P� �;6xy�u�z�7jd���	��uuL5U�P����G���Scd�yc�E��VY<Fx����ќ�-��#���0/V6#V:�܆�I>f�o)������zO�xL�� ���fttȪZheO���j�0b=p��.dgKce���'���nOv�EQ�9}�&�Q|X��� �y�K]5�X�5ʃ�F��1C49H�j� �͍�$~���HoF� VP%}��d��C�c<�}��@� �#'(����~��r~Ei�aqf���<�+�N���X�[��D5���4}Y��ft��GR���r���OtB��Sb|�x�Z�u�����)�U��6)*PR�%`��k���^�����K�q�Yd)d(fФ)en2�ImX�s�Ʊ��H�����!߭T�P���'�(�x*�����&�b��=� ?���?}cb
��;�D�go���,��r(C;�r1�z�v&�'}��J��!xI!��ms�K���9w�տ3�3�t�w�"-����� �v�J��h1�v��t]t4�'Z�:C!9NX���,B۰Y�W(�/,K��gF�4I$�<[�q��U�뱡7=����<�pX�Q��Eb�MJ�@ )142�䤋
�n���J53�/$�DU6���C�Ҽs��}-;P]zg��j��A4�M��{[������D����R�n�C(<g��G�k��uүä�	�V��%�9]w�9��.r$��P3ۦ;�֌$Hk��j�49,�Z�}A{d��/H0rV�h����TA�e�S��4��m9i,K�K�#���,��3�>� )�3B��d���Zc����[CD_`n1�Rңo������$��"[�� l��{i�&�%(�J����z�A���Aj�2x�ao�^T����m�˺��R��8��ǭv�����l蒚�jlMv*ĸ�8d&�U5�$8�����Ԫ]�G�D��#��l��(&/I���5h�X �ܵ��!6pR0v�.|l},�J��e����w�6�n�M9̔�Ahq��G׺V�K�������_��[6c��G���
�[��Ǚ��Zl�;�>��9�ԛ
���REfh�]�g,"A�1Ku��l5
��撉ي�,�.9��L�T����B�B����vk]4�%&3��L�hoK�Ƶ�`|v��_�.���j���Fk��W���8Ӑ;��Ck����a���E�ĳ�
}<�\��'�qM=���܆0
���^�8%�+[ !�vX�`C.�N�E���������!~�s��_?�7��\:ܔ�pG\�5W��MBA��ѻ������\ِ�5w�APX�ͧ���o��5JW��^�0 ��AM�5�h	�	�cFVw2U���yug��:���Qa�:`f�y�r��?��#6?����I<۩��Q��K:H����!�'ޜj�h~�O����^a�4�̽]M��ӆ���wy������Mc�S;o�.
����{�������w��͢��q�G�dɆ��b!�0<���sR|��1�B��3{x�>=$,�H.���R;��
��w3���J��w\��:x�*��^h���ni~r4T*�'�z���T�*������Zl|6䱗��r��;����q��r4��f��\��V�9Q�)��|x������2��$dUL�!k'��ZT������7����-xݯ��������ϐz\N{R�� h�߆�jun.ښ7�&���y���4����ti�7+BX�4�u�+nv�p�V\g�7)e7%g�1�Ҷ�'7��<���5�{�����u5%���ݵ^a���1�H/�Z1ď��y���>G`�y�\���D��asE�(c� ������ηlK�z�S�զ0�yB���
���5�M�^�������a��ׄ��FdWM9(��Gj�H�$������:n����$c���e\O�G��eTX[×�����]Z��
������X���H "3��Y?��q+zĢ]_�3�ڸ�"aoU��Eā��Á 1�:���������k�w9/�qE�HRzbtN�x�F���6Z4��v�wԺ���_�>�@���b�1e�+�q����+X�Z�[�+��cp �D�)k�m�CS>�Zq�3�ɶ��I�im�dE�_ݚ�d�pk6�L��r>k��O���x?� �{nk���[m�85��!������f�I�~d�º��aV���nuΝ��/c/3Fc-
�9��q���<���`�(ewf�LY �UBm��+},����K�)��	��"	��<��H�-��:�z��/�}qlˊS�������L��$P���Kc
'��ƨK�"�>��ɢG�R-9GP�$0��]�Ik�h1�����(ޅ<�>Ck$��!�+HN�B|����L�M�IY���H(m�?�&II��J�� ͋F`�������*��*��l ޼�"�3[��"��L�=SZ@!�=�Θ41��c���ĜvE�;D�N�����J��1�(f�Υ�y�_z����I�F1Q^[4���t�$�,�������dR�qk�9�k-�W�HD@�
�&���^o���n�@�w�L��ŝ@�#����ƃ�������B ���{L��:�5�����oPHg��J-������F������i
ڭ��Iz�]Ar�^�bm{ H�l�d���Q/y�&�<U{���)ɇ��	��p���J⡾&��iAk0��R᫣@����J#��>��R�8&Q	�?�ݨ�l�"����dlޤ@�&������@� } ��7��+R�¾2\�G���Tf�Y���q������oV����SڱHgvw#vw��J���ȧ�<'RB1� ��4���Ouw��./$����mIT�H{���d	�a�Z�V9��_�d�quV�~H���-ʏH�� �d,�:e̫��u��$S�� t.�,f�	ї�'��l�@��8����ȍwEGⓞ����T:�p?TL������K �%Ϭ7�Q|��HGB��z��H�m ۙ��<�����$��s^}x�O��Zn�?�'��O4N��n�=�c�����H�Ǫ��[�t0`�h��`^h���k��<��2�,�h�b�9��V�M�f�*/��ZԼv�tFk�ܱv=9��J�| /+q�.��(��Fy5ؐ:��h�a�kBOc��n�^�hh��������������l'B�t�H�~Z�+�XZ���$��xf!*H�q��b�$;��3nXZE�W}�p��ݠ�˃N�K��X	����J�-�l�W��_+�^`m��7����-��J�Z�/�81�Ի�m�
	g����q��� �y�����(��b�Ky+!�T#�W} �5�13)�q/�f�L�N"��o�|�k5ـ�X4[ �>8f�am��S9e[j��E4��:}���<��X�ű,s!�<ҢP��6��loБ��d?R��j4m�{~N����(�d �����N�F@!��0��S��Ѭ�|WyX�ڐ/��k��=��s �@��ć?GPE�x�ȴB8>�G���� Y/�gLD�M$�Hβucg#v7���:̶���4���>�ޔ<]��?w�N���F�?�)�_�`���哾�����Az�ɉY�u�}H��#�yv�+o�:kI�������x����~��}L�d�G����1끖��d�I�@�B+�g��(-�П`|��l�o�C�_�B��yYΦ[C�A<��2���c}
���ő��K��,���f&+������Z��<�Й����N�����m��)p\�>�T ��qP���Mא��"� s���"�u���}�+߮�qV��Pެ^��t���W�c���8(����&(�+���M�O�n��I��@N,�]#m���xب��N&k�[�����E�o��r���]X�e.$���0)f>�������c�ɐ����R���I>*D] �*T�a]�O���8L=��ؗ؜��-�,�5�slc���&��!MSbr�$����q/�_X�>��PQo��AƷvm�L�00Y���P� �� ��M"L�ǎ��)����|X�n�i�0�Oa�/8�����~�b I�w2�)���>�B���.e۝����X�W��	�䥛�xmv�+�u�M��(j;"�͗N���\�Q������Y�@�)�{�I+��0��P��q�Q��M��2�����`��j��W%r��`�������۵x5ӖE!]����1���ĶO�oD�Ҋ%N�Yf>��`Qcz��$��ea��	�y�Lc�W@'3Mi���Ul�9\F�t����uظ��Hv�myA�kcQ�����j,<R�k����btbp�� ��\���f,[�Uj��c�a�]4tGx�~TA#�G���5�'�ҷ�&w[�*��{�˃]����*�����7�4;5���>�Uij��i���X�=��D�����-��X"$�Rovv���I�ɮ�"L�E�Mͯ)|!�Hw	(��P"ӃT�yIn�82�Q��}�.%Ŋ�_��f�Y�/�(�4	m��,I�W1�YHV�?��Bx.� ��_��rI����јn�yCCvy�)�3 $��`��1[�� ș��h�A�~b������7�I�����
��{��Y�3�8��e�
BOf��O�u�;~�C�Tb+���mB�M���B��KL\Kw�e 8��G� E�sഓ��qA��a��� W����z�?�eJ	��kw�����g!{u�`���\e�y���dz0�?�Aـ�'yd;-�M����f f�=\�q���"�uI"23L��ϑ9� P*���}q?'��V�u0i��LQ˽�S#�`�p_5d�@;_��x��0.Ff#���N��(Al�ۘҁ7ʏ!
5�+B[����E2�8��N�$�!��Gt#����]
4�l��NN�qc�����-���?&�L����<v��*������NF>>B�b�O����F}��~��1�5�61]�EI��CY�w��������`��z ���S�����p�I2�VHe�oc)5��'�d07-4�5I�@��i!b��h`^��i�w��V�˶j�9D�K�x����J�L��}���p���z��L�0;�}�҈0��L�%���\��ͽ�� �a_�Eau/m�N�r���Q�0����Zy��D�.l�$vT���� �닢:���~�Ⳅ�\�b��#�Ʉz�%�2܈T]��n�cz6�R|�E��49H�ܒ��a%h�oƝ���_��&�&�8�"*�慅��A�P8�ச��T�I�X���?�9����2A������v�a�$�K�������
��h������l�\����*h߅��c��c�����I ����tf6�<JL$-�?Ϣ�,4S�!�1NJ�k$v�s��;��.�'�kmeb�T��V��,Xچr���oO��	>>墏�+e�<������R1��l���c{94CbI���Z������7��Z�6��&�҅ٞ�`T�a�V$x~��V����+T����v�}����C�mj�O8d$���63�&%�)=��t
P��{�@8^c�)E0~��t���lL���ɻ�I���=���֞����>�K�_�d���d�+Ey�	?�nhc���L&�ݟYH�N�%�d�+U�
��� �\2�54�x;���G�2�&�~�� ���ˑy��UN�f5���r`����'��c��C�W����!�/�J��C�sJ��}Z%�����T�e��(�vP1.kC�^MM"��nQh��d���,�ZD��t�))G={�����2�.�q��GMm*ҍG�D�������xV�p}�ʎ>�`B9Y�r8��T�蔚uI�Nw�UVu���J@v�8��9�WRL��Ci}�
�m����v��aG
�p��'
��mR��ư�N�:��Z�J�����Vc�֝��aU�$�6��h�
��ح�_�
��
�����_������� ~5�u���^e�|E�N��f����Ug^�� %�~���%fTӅ��z@�b�2ɞ3����u����ŉ��	��Z��!W�C��a@zn����@�l\� �p`?��5B��K�>\�kEٶ><ݧ�0�qm�k������E�\�����!F@�yw���� �'��y/��[2��
"Mnn�X7�:)HL�o&�j:�f#���.du�;\�z���9����y=��s�_ZP�G半�	���\L��食o؍��QipU�?_a�S�;{���C���:
cI��U��k�#ʝĚC��`���F�Wg��?�t삕v�25�ub��+d�=&/�fQ3�~U�NMadj?@�~��I�x!����%�«0�Z�ÛD���A<ٺ�*`��a!��vռ1RV�B��|c`��b@f�y�[�Fk��C(#\�`!��'܋�Y�Ca�&�ʎ����V�n�j7�9��������~���"D�<Ν��T���^��O������7=^G�����S=�K�����x}R�4{<��W�{�N���	Uv���^n����������;�C�j�Kz;}����~�'u��?����ƦB�,!M˯����63��d�W[�~�]���$s�	��y�"[Q�F;+�Ev�����,&qع��frDs�������X��[9TSi�_s��;�t�o�d�~�O]Meb�:�d���������͕��v��%�{�|�)���)��]2���/?�_ʦk3$�k��P�s�ʚ�fms_�Q;+�Xy.�
���t)Z�&U--̎4F�:�_J�yD��-�Ђ/���X�z���i�Q<�#��S��;�3r�$*���w�g�Ԟ�>g�]`�p�[��: !�6�G��?;�$�j U)*��4Wl�b��� -��X�&����H�0����Y]{L�;k��V��oC���lcdv����-�ZA6]���Q�q�l��^�V(y��mq���AW�Q�Sލ5� �AM��	�qMr���Y0{<�r���Lx�ڂ���^6j& ��A�Y*��-��P7�M���x��R&��D {�S����F�^��p�S$.�'!��n�߇A��TO���V3�?�(�,8�����"��'8������p���t?�T;
�����Sh3��+8��DTdJL��"��?ܟ�+t�DFo��=e"Ч\Q��72�f�������!�ݫ�nm.�Ѯ�ŮC��)	>�Ӌf+�эmu����3���`�+^t�;O%�HQ<l&)�,��Jo��F� ^�Y�7tF�!�}l���-0ؠ~s�<�iF#m겅�70��u)����\�/��<���P�����?��q��b'?K���x�d���B2o�z�^��q�E;�f3x��� b���*�f�=��on9��>?����L�b�X:�AB�w#��Dٌ����7�Hpqvq��2���&��8Y�#��������S�u��"����7� `Z&F7T�XTX�*p��R����|�48�|D��Bg�f,D��1y̩-S[0�?JW�X��"WC:��w��|t�R�?�<�(+㘁K���h?�K$�/�>�%�f�te��Fh���s�N*��݉�AhB/#�31���=�	�;�`J4�}��g��H���u����w�C�䭟����.���kG����Z�/�;rs��w*NG�e�m-|��c�ԟh�|t�R�J�o��l�nc��	�A���_�� �}��<��V���P����Ul}|/�{��x�e�$e	+��`�߉￶;����b�g5T����z�����zx�����	���_��hr6�Gi�,P��P@y.@�ԟ����.��y�-4��/ζ�!�W��,[^���p�@l�}Lm6�n Y�*ʠ���j��q�zG�k;k���tn��A'��=Қ=F%��u��V!q�*��t�c�N�V�V7̶�*������u��y������`�J��3����Xʞ�ŋ����?�U������}*F<���՚ruY�R���2HGC��s�����sa�:d�޾TX��Y(��RT�:�!mo��ݙ����i�1�W��Ժ�k�z�qL2�۪,�Y���3ާ�e��
���'X�����r H����_�Zop�g��0�����|�#FD��Z��8�;� vϑ{{�tW�핆��`�����8k�h���i��qS#΁Pc$�VP��HuwɼDL�<��jM�ҽ���J�O�k�~ ��z=L����O�����?�0�T~���+C�.5z�/��t�a�,F<~��L�ݕ��H�$W�P���g�g94K���ϲ<��j�|I�u�I�A5�#�Z�XY�D*(�� ���2�6d����\���;��8���m`�����gf�/� �l�Y1��9�ш>��b^�T�5������"t}���ql��K&�e�8��3Py�RӣX����c��1�*��gũ�D߻�lbE������(�k@2������=EE3�����۔w ����~"%��r�wi�!#;U.�l������CDJMX9VH�`�J���M�ӡ�r�Dl���wT4ŋ`��(D�?	z'�^�)�t
����^R��˟�9W���c�2�B�����b��7�P��r��S���ئ;7�`�ŶK��#Z(^�ȷ�������%��o�ϗV�����M�W�	�/;Q�)�8"�Ca_�!�'���K�;<�Q"��u2���6�nw����;���.>��8�r5��K3a��&��p�8n��,T�G5�s�q���3��0���f�Z�qG��'�{�3�tu�)���HQ����'����
�X&1����E�}־�wj�g�����d��(���AɄF�=� ��j��*l�@J��S��o�b[ �`籿�ZR)������{@6~�V�b1��ϳ6�ĤK�����8��h2�l#F�H��G#GCZ��ͳ!X���V�
5c�~�ҲE2A�����dE�.�W�\�=����!�%3n�b< �?`r.�OWB��|O�qzwC�6�~u�03�z)XB������؝�Zƚ�#��uϩV`[o�2!�m�v��+�	�i��`|��3��f"|M~��.RU�p�mQ�?��̙�?ϙU
T�!E�ÿ`|)ݸz�d߰J�9�^o�{q�U
��N�U�GֲJ�����Ww��jB/ė;�fM�nL%�U��B'�"�F�и�ᥒg���c�IN��	9��CǠ��؋%�q�ލl	O�Jaf�Sl�d����49P-^�=��$��sb�c�b�s���e���;��&�����&��v���Ӻ����L��$~ς�+r���j������ڽ/VdN!��j���Q���c�2�����"�����6��.&NW�Xc�D�"����W�?���Y@hy `����"�ô]�T,�+ے9�u@!��>�~�D���c����F�X�h&Z�� ֽך(�L�-k�&� 9[ů2�zUK��Rc��<�mi`�&Q�
�!�3��	�ԏM��4m�w+�$9�rY�oF��qա����)�|�^�g�a�B9��E�0�����L5�����Alpx޸$ٰ�ѥ��0����b_�lCM�M���Ƽ{���<V��gk?�W�5����Bg����ԩ��B�2� lm8�B���Ӈ[�$_=�X�Ş�:~�ܠ�g+�^�C���|�$4c#�F�Qw�]�oj�6u۹T�O��l�o�G��x����������m fv!�ִ����vE�}�NLG�;�ȕ-�G��t���
���Ƴ�L�̦:�j1�����W��,`���?n�XߎC�s��r�L8�"Unj��x�IkS|�� NocCG��}�����R*#CTD��F�\����6�w�����2��#`5iB�r����<���(���dG��~���VK��k�L6N(dQ
�'ٶ�{�2<>���|��#ڻ(���h1S=�64�ӱ��?�)�Hi����B�A���]����5�B���ޱ+�WnX���2��F���h0�S��t½�%�����#W�*�
j�)�x��8�}���A�'������nv'�n���e�qI�A	��.�U�ɰ�k�2o�t�$/���$�1	�릙�լ9�qt��(����"l��~*h��wo*��%�]n�xW/��� ���ʫ��v*#�3��:��&3��k������"����D�|f���[�O#b�0��Ƶ�ݹDxT6������\;s&}���.��iu���#�����ˢ���z}�\�E��8�|�=��B�%����?;�G =�u��:��ށ:������{���P���J�� |��o���,dҀ��sC~h��)<�c*�%*л}`Z�_�0EM����0I���6]Z��3������A����0v��2d�.�|R,��ӟxFt��,�t�m��;��K]��������>�{ch��0+/Fh>Ud��?s�����w+��7=�d�۟�'��6�p�c��P5��k��.����K�c��g�9v�a�p���n&�E�7A�iq�Zo�Zas���[��>̕�[+��
���Y�N��E�0���ma]�c.)���:���S'��5�RG�癤��SQ�S�<U��	9
��S�>��/V��J��?a�wx��ɤ`\�Bڳ�7^���$h.�6��w��̑E�HYiQ�����bٜ��	�~1�٩���H@����������3�+Nw��e��,M�Dvcl�v^����fi��_!�����-�k��
�4.g�^���R�Sϋ�f��G����۫]�?��.��w-׌��i�q �y^�����1�>_��� ŦBpV�<��y�,�֑�����v����9`�>�ҎH:��f�:"�uŤ��k~G� ~�9�,�<5�0�:8�4�]0L�[.zm]��Me�U��vaЯ�5$��>�,f�#@E޸�:��rń�F��Վ!�����\2��FiA�`�3��z�l����D�'��p�|z����ڃk��S�N(�yp��\��f�
�>�ʿ�6m�7�l1���)YGV�u�w�;�g�r5;�K��/N�i3�7���b	#��rr��*���Б�y(�����pu�,�)����y���_-��fq���YWފ�&��A(�阔����1���e��I�z���^�4��>�g��ɞ��
n�i����(�^a{v�Y�g2��pb&�"K�j�^>��m��.�=j��x$�)�M�QEKs�
t��p�Q����YTe	�u�ʜ�=�j��j�(w����/�0 :��h�����@G NЌzsb�Q�.Y�����
0'(��ה!�(6o\������r(6�{�xr�(ߐI��V1 JU�E��:g~-��<٨��m��C�M�2�D*�D����	���K~vj�r	�rv��V�-��CR	��E���H6mN��նL�$�G!l��ӅR�Ñ}ꢕ�ó�LGS�w笒��������^��-����ՎTc|���IoJ��ҩ�hm�_�7
��^7!�_,�R��ԯS����+�y�i�ht@�.YC;�K�ԭ��4�����Q!��Z�.�}�v�O��/S�{0�&p�س��)�RA��dGJ�b�	��3�r!"$�,|�9Q�1�^�}�M�C<,{<��Q�h�4�.�Y��O�D�}��$`:p��>/�Ъ�S��%q��>�m<��{t6�#S!��؈�𼶑J�H��aA��� k�@P��0��uB����g����h�ԑ�Q����t���m�"�+ur�_ӡ�=frM����u�Rp�TZo�����ʆ����4�cr�2��桔���E�<���2rI_e�G��[ x��eFz��Q��2�+pk?Bi]D|�5C;ORtz�tu��(�6'j"�<��A������r��;����h"x*��%�CL���S�8�Aj����l""ae���H�֑�gو�i��ٿ���(_y��-q�Tf�jOUen۱�g��E��N
���K�^��<@�x
�=�ؘo2�Nli�&{NZ�o��"�_q_����P6��w9D��
������S)'�/�B��w5y�`3���j�x��oh��˛V��F]�WP�Э��?���~Kj���F��bu���d�<����H�/7�&|�3N�g�f�)�۵s�O{Z���V!���\��;�ѱ�s���ɞ����B�6���G;��o��� Y�G��iT�0���_#�;�?����%Z�b���ʖ>�,���J��g&�&'6c���;��apEK���	���*�+������].5�Ö:^\87y�f<��p�X�#��񊣄[����$l[��6;i�,@��
��"�	���#�6�+$!�Ә�Q�P�D�=f&L�>�_S�(d�/��w��K��*�Ow"+]�)��
����A���B�og�:=�L��j7axe���0���>]1��J@����r���%��ӝ܉9-�uy��8�3�ê�Z]�쿗�m`�J1���_����
�X11���$���'��<��~�oWaV���kl��Û���o�/<�39'�(���<O�V�h���P��q���*����ޝQ��&�JK��rl���3Y���U��>KVO v��<�FZ_|��g����ȡ���_��:���~���n͇^��T�P�XZ���C�ōO)�&Uc=�n^�aE��0����q�����M��x�c�B/��� �6���&AgB'"&��m�^�Z�]/ �J,����W��H/�M�Y�F;(��(G14��Eӆ�rW鮴s�	ƌ����?��PPyZf?'aW�0I��r,z?1��}��c����B( ��5~�[�\$wu�\K�'���A����O�N�4p�ӎ�2V��uTA|ueX���jM�׊�
s