// deca_vip.v

// Generated using ACDS version 15.0 145

`timescale 1 ps / 1 ps
module deca_vip (
		output wire        altpll_mipi_clk_clk,                           //                 altpll_mipi_clk.clk
		output wire        altpll_sys_hdmi_clk,                           //                 altpll_sys_hdmi.clk
		input  wire        clk_clk,                                       //                             clk.clk
		output wire        clock_bridge_vip_out_clk_clk,                  //        clock_bridge_vip_out_clk.clk
		input  wire [3:0]  ddr3_status_external_connection_export,        // ddr3_status_external_connection.export
		input  wire        hdmi_cvo_vid_clk,                              //                        hdmi_cvo.vid_clk
		output wire [23:0] hdmi_cvo_vid_data,                             //                                .vid_data
		output wire        hdmi_cvo_underflow,                            //                                .underflow
		output wire        hdmi_cvo_vid_datavalid,                        //                                .vid_datavalid
		output wire        hdmi_cvo_vid_v_sync,                           //                                .vid_v_sync
		output wire        hdmi_cvo_vid_h_sync,                           //                                .vid_h_sync
		output wire        hdmi_cvo_vid_f,                                //                                .vid_f
		output wire        hdmi_cvo_vid_h,                                //                                .vid_h
		output wire        hdmi_cvo_vid_v,                                //                                .vid_v
		output wire [7:0]  led_external_connection_export,                //         led_external_connection.export
		input  wire        mem_if_ddr3_emif_pll_ref_clk_clk,              //    mem_if_ddr3_emif_pll_ref_clk.clk
		output wire        mem_if_ddr3_emif_pll_sharing_pll_mem_clk,      //    mem_if_ddr3_emif_pll_sharing.pll_mem_clk
		output wire        mem_if_ddr3_emif_pll_sharing_pll_write_clk,    //                                .pll_write_clk
		output wire        mem_if_ddr3_emif_pll_sharing_pll_locked,       //                                .pll_locked
		output wire        mem_if_ddr3_emif_pll_sharing_pll_capture0_clk, //                                .pll_capture0_clk
		output wire        mem_if_ddr3_emif_pll_sharing_pll_capture1_clk, //                                .pll_capture1_clk
		output wire        mem_if_ddr3_emif_status_local_init_done,       //         mem_if_ddr3_emif_status.local_init_done
		output wire        mem_if_ddr3_emif_status_local_cal_success,     //                                .local_cal_success
		output wire        mem_if_ddr3_emif_status_local_cal_fail,        //                                .local_cal_fail
		output wire [14:0] memory_mem_a,                                  //                          memory.mem_a
		output wire [2:0]  memory_mem_ba,                                 //                                .mem_ba
		inout  wire [0:0]  memory_mem_ck,                                 //                                .mem_ck
		inout  wire [0:0]  memory_mem_ck_n,                               //                                .mem_ck_n
		output wire [0:0]  memory_mem_cke,                                //                                .mem_cke
		output wire [0:0]  memory_mem_cs_n,                               //                                .mem_cs_n
		output wire [1:0]  memory_mem_dm,                                 //                                .mem_dm
		output wire [0:0]  memory_mem_ras_n,                              //                                .mem_ras_n
		output wire [0:0]  memory_mem_cas_n,                              //                                .mem_cas_n
		output wire [0:0]  memory_mem_we_n,                               //                                .mem_we_n
		output wire        memory_mem_reset_n,                            //                                .mem_reset_n
		inout  wire [15:0] memory_mem_dq,                                 //                                .mem_dq
		inout  wire [1:0]  memory_mem_dqs,                                //                                .mem_dqs
		inout  wire [1:0]  memory_mem_dqs_n,                              //                                .mem_dqs_n
		output wire [0:0]  memory_mem_odt,                                //                                .mem_odt
		input  wire        reset_reset_n,                                 //                           reset.reset_n
		input  wire [1:0]  sw_external_connection_export                  //          sw_external_connection.export
	);

	wire          alt_vip_vfr_1_avalon_streaming_source_valid;               // alt_vip_vfr_1:dout_valid -> alt_vip_cpr_1:din0_valid
	wire   [31:0] alt_vip_vfr_1_avalon_streaming_source_data;                // alt_vip_vfr_1:dout_data -> alt_vip_cpr_1:din0_data
	wire          alt_vip_vfr_1_avalon_streaming_source_ready;               // alt_vip_cpr_1:din0_ready -> alt_vip_vfr_1:dout_ready
	wire          alt_vip_vfr_1_avalon_streaming_source_startofpacket;       // alt_vip_vfr_1:dout_startofpacket -> alt_vip_cpr_1:din0_startofpacket
	wire          alt_vip_vfr_1_avalon_streaming_source_endofpacket;         // alt_vip_vfr_1:dout_endofpacket -> alt_vip_cpr_1:din0_endofpacket
	wire          alt_vip_cpr_1_dout0_valid;                                 // alt_vip_cpr_1:dout0_valid -> hdmi_cvo:din_valid
	wire   [23:0] alt_vip_cpr_1_dout0_data;                                  // alt_vip_cpr_1:dout0_data -> hdmi_cvo:din_data
	wire          alt_vip_cpr_1_dout0_ready;                                 // hdmi_cvo:din_ready -> alt_vip_cpr_1:dout0_ready
	wire          alt_vip_cpr_1_dout0_startofpacket;                         // alt_vip_cpr_1:dout0_startofpacket -> hdmi_cvo:din_startofpacket
	wire          alt_vip_cpr_1_dout0_endofpacket;                           // alt_vip_cpr_1:dout0_endofpacket -> hdmi_cvo:din_endofpacket
	wire          altpll_sys_c1_clk;                                         // altpll_sys:c1 -> [alt_vip_cpr_1:clock, alt_vip_vfr_1:clock, alt_vip_vfr_1:master_clock, hdmi_cvo:main_clock_clk, irq_synchronizer:receiver_clk, irq_synchronizer_001:receiver_clk, mm_interconnect_0:altpll_sys_c1_clk, rst_controller:clk, rst_controller_001:clk, rst_controller_003:clk]
	wire          nios2_gen2_debug_reset_request_reset;                      // nios2_gen2:debug_reset_request -> [ddr3_status:reset_n, mem_if_ddr3_emif:global_reset_n, mem_if_ddr3_emif:soft_reset_n, mm_interconnect_0:ddr3_status_reset_reset_bridge_in_reset_reset, rst_controller:reset_in0, rst_controller_003:reset_in1, rst_controller_005:reset_in0, rst_controller_006:reset_in1, rst_controller_007:reset_in0]
	wire  [255:0] alt_vip_vfr_1_avalon_master_readdata;                      // mm_interconnect_0:alt_vip_vfr_1_avalon_master_readdata -> alt_vip_vfr_1:master_readdata
	wire          alt_vip_vfr_1_avalon_master_waitrequest;                   // mm_interconnect_0:alt_vip_vfr_1_avalon_master_waitrequest -> alt_vip_vfr_1:master_waitrequest
	wire   [31:0] alt_vip_vfr_1_avalon_master_address;                       // alt_vip_vfr_1:master_address -> mm_interconnect_0:alt_vip_vfr_1_avalon_master_address
	wire          alt_vip_vfr_1_avalon_master_read;                          // alt_vip_vfr_1:master_read -> mm_interconnect_0:alt_vip_vfr_1_avalon_master_read
	wire          alt_vip_vfr_1_avalon_master_readdatavalid;                 // mm_interconnect_0:alt_vip_vfr_1_avalon_master_readdatavalid -> alt_vip_vfr_1:master_readdatavalid
	wire    [5:0] alt_vip_vfr_1_avalon_master_burstcount;                    // alt_vip_vfr_1:master_burstcount -> mm_interconnect_0:alt_vip_vfr_1_avalon_master_burstcount
	wire   [31:0] nios2_gen2_data_master_readdata;                           // mm_interconnect_0:nios2_gen2_data_master_readdata -> nios2_gen2:d_readdata
	wire          nios2_gen2_data_master_waitrequest;                        // mm_interconnect_0:nios2_gen2_data_master_waitrequest -> nios2_gen2:d_waitrequest
	wire          nios2_gen2_data_master_debugaccess;                        // nios2_gen2:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_gen2_data_master_debugaccess
	wire   [30:0] nios2_gen2_data_master_address;                            // nios2_gen2:d_address -> mm_interconnect_0:nios2_gen2_data_master_address
	wire    [3:0] nios2_gen2_data_master_byteenable;                         // nios2_gen2:d_byteenable -> mm_interconnect_0:nios2_gen2_data_master_byteenable
	wire          nios2_gen2_data_master_read;                               // nios2_gen2:d_read -> mm_interconnect_0:nios2_gen2_data_master_read
	wire          nios2_gen2_data_master_readdatavalid;                      // mm_interconnect_0:nios2_gen2_data_master_readdatavalid -> nios2_gen2:d_readdatavalid
	wire          nios2_gen2_data_master_write;                              // nios2_gen2:d_write -> mm_interconnect_0:nios2_gen2_data_master_write
	wire   [31:0] nios2_gen2_data_master_writedata;                          // nios2_gen2:d_writedata -> mm_interconnect_0:nios2_gen2_data_master_writedata
	wire   [31:0] nios2_gen2_instruction_master_readdata;                    // mm_interconnect_0:nios2_gen2_instruction_master_readdata -> nios2_gen2:i_readdata
	wire          nios2_gen2_instruction_master_waitrequest;                 // mm_interconnect_0:nios2_gen2_instruction_master_waitrequest -> nios2_gen2:i_waitrequest
	wire   [30:0] nios2_gen2_instruction_master_address;                     // nios2_gen2:i_address -> mm_interconnect_0:nios2_gen2_instruction_master_address
	wire          nios2_gen2_instruction_master_read;                        // nios2_gen2:i_read -> mm_interconnect_0:nios2_gen2_instruction_master_read
	wire          nios2_gen2_instruction_master_readdatavalid;               // mm_interconnect_0:nios2_gen2_instruction_master_readdatavalid -> nios2_gen2:i_readdatavalid
	wire          mm_interconnect_0_mem_if_ddr3_emif_avl_beginbursttransfer; // mm_interconnect_0:mem_if_ddr3_emif_avl_beginbursttransfer -> mem_if_ddr3_emif:avl_burstbegin
	wire   [63:0] mm_interconnect_0_mem_if_ddr3_emif_avl_readdata;           // mem_if_ddr3_emif:avl_rdata -> mm_interconnect_0:mem_if_ddr3_emif_avl_readdata
	wire          mm_interconnect_0_mem_if_ddr3_emif_avl_waitrequest;        // mem_if_ddr3_emif:avl_ready -> mm_interconnect_0:mem_if_ddr3_emif_avl_waitrequest
	wire   [25:0] mm_interconnect_0_mem_if_ddr3_emif_avl_address;            // mm_interconnect_0:mem_if_ddr3_emif_avl_address -> mem_if_ddr3_emif:avl_addr
	wire          mm_interconnect_0_mem_if_ddr3_emif_avl_read;               // mm_interconnect_0:mem_if_ddr3_emif_avl_read -> mem_if_ddr3_emif:avl_read_req
	wire    [7:0] mm_interconnect_0_mem_if_ddr3_emif_avl_byteenable;         // mm_interconnect_0:mem_if_ddr3_emif_avl_byteenable -> mem_if_ddr3_emif:avl_be
	wire          mm_interconnect_0_mem_if_ddr3_emif_avl_readdatavalid;      // mem_if_ddr3_emif:avl_rdata_valid -> mm_interconnect_0:mem_if_ddr3_emif_avl_readdatavalid
	wire          mm_interconnect_0_mem_if_ddr3_emif_avl_write;              // mm_interconnect_0:mem_if_ddr3_emif_avl_write -> mem_if_ddr3_emif:avl_write_req
	wire   [63:0] mm_interconnect_0_mem_if_ddr3_emif_avl_writedata;          // mm_interconnect_0:mem_if_ddr3_emif_avl_writedata -> mem_if_ddr3_emif:avl_wdata
	wire    [2:0] mm_interconnect_0_mem_if_ddr3_emif_avl_burstcount;         // mm_interconnect_0:mem_if_ddr3_emif_avl_burstcount -> mem_if_ddr3_emif:avl_size
	wire          mem_if_ddr3_emif_afi_clk_clk;                              // mem_if_ddr3_emif:afi_clk -> [mm_interconnect_0:mem_if_ddr3_emif_afi_clk_clk, rst_controller_007:clk]
	wire   [31:0] mm_interconnect_0_nios2_gen2_debug_mem_slave_readdata;     // nios2_gen2:debug_mem_slave_readdata -> mm_interconnect_0:nios2_gen2_debug_mem_slave_readdata
	wire          mm_interconnect_0_nios2_gen2_debug_mem_slave_waitrequest;  // nios2_gen2:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_gen2_debug_mem_slave_waitrequest
	wire          mm_interconnect_0_nios2_gen2_debug_mem_slave_debugaccess;  // mm_interconnect_0:nios2_gen2_debug_mem_slave_debugaccess -> nios2_gen2:debug_mem_slave_debugaccess
	wire    [8:0] mm_interconnect_0_nios2_gen2_debug_mem_slave_address;      // mm_interconnect_0:nios2_gen2_debug_mem_slave_address -> nios2_gen2:debug_mem_slave_address
	wire          mm_interconnect_0_nios2_gen2_debug_mem_slave_read;         // mm_interconnect_0:nios2_gen2_debug_mem_slave_read -> nios2_gen2:debug_mem_slave_read
	wire    [3:0] mm_interconnect_0_nios2_gen2_debug_mem_slave_byteenable;   // mm_interconnect_0:nios2_gen2_debug_mem_slave_byteenable -> nios2_gen2:debug_mem_slave_byteenable
	wire          mm_interconnect_0_nios2_gen2_debug_mem_slave_write;        // mm_interconnect_0:nios2_gen2_debug_mem_slave_write -> nios2_gen2:debug_mem_slave_write
	wire   [31:0] mm_interconnect_0_nios2_gen2_debug_mem_slave_writedata;    // mm_interconnect_0:nios2_gen2_debug_mem_slave_writedata -> nios2_gen2:debug_mem_slave_writedata
	wire          mm_interconnect_0_onchip_memory2_s1_chipselect;            // mm_interconnect_0:onchip_memory2_s1_chipselect -> onchip_memory2:chipselect
	wire   [31:0] mm_interconnect_0_onchip_memory2_s1_readdata;              // onchip_memory2:readdata -> mm_interconnect_0:onchip_memory2_s1_readdata
	wire   [14:0] mm_interconnect_0_onchip_memory2_s1_address;               // mm_interconnect_0:onchip_memory2_s1_address -> onchip_memory2:address
	wire    [3:0] mm_interconnect_0_onchip_memory2_s1_byteenable;            // mm_interconnect_0:onchip_memory2_s1_byteenable -> onchip_memory2:byteenable
	wire          mm_interconnect_0_onchip_memory2_s1_write;                 // mm_interconnect_0:onchip_memory2_s1_write -> onchip_memory2:write
	wire   [31:0] mm_interconnect_0_onchip_memory2_s1_writedata;             // mm_interconnect_0:onchip_memory2_s1_writedata -> onchip_memory2:writedata
	wire          mm_interconnect_0_onchip_memory2_s1_clken;                 // mm_interconnect_0:onchip_memory2_s1_clken -> onchip_memory2:clken
	wire          mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect;  // mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	wire   [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata;    // jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	wire          mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest; // jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	wire    [0:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_address;     // mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	wire          mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;        // mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> jtag_uart:av_read_n
	wire          mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;       // mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> jtag_uart:av_write_n
	wire   [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata;   // mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	wire   [31:0] mm_interconnect_0_alt_vip_vfr_1_avalon_slave_readdata;     // alt_vip_vfr_1:slave_readdata -> mm_interconnect_0:alt_vip_vfr_1_avalon_slave_readdata
	wire    [4:0] mm_interconnect_0_alt_vip_vfr_1_avalon_slave_address;      // mm_interconnect_0:alt_vip_vfr_1_avalon_slave_address -> alt_vip_vfr_1:slave_address
	wire          mm_interconnect_0_alt_vip_vfr_1_avalon_slave_read;         // mm_interconnect_0:alt_vip_vfr_1_avalon_slave_read -> alt_vip_vfr_1:slave_read
	wire          mm_interconnect_0_alt_vip_vfr_1_avalon_slave_write;        // mm_interconnect_0:alt_vip_vfr_1_avalon_slave_write -> alt_vip_vfr_1:slave_write
	wire   [31:0] mm_interconnect_0_alt_vip_vfr_1_avalon_slave_writedata;    // mm_interconnect_0:alt_vip_vfr_1_avalon_slave_writedata -> alt_vip_vfr_1:slave_writedata
	wire   [31:0] mm_interconnect_0_sysid_qsys_control_slave_readdata;       // sysid_qsys:readdata -> mm_interconnect_0:sysid_qsys_control_slave_readdata
	wire    [0:0] mm_interconnect_0_sysid_qsys_control_slave_address;        // mm_interconnect_0:sysid_qsys_control_slave_address -> sysid_qsys:address
	wire   [31:0] mm_interconnect_0_altpll_mipi_pll_slave_readdata;          // altpll_mipi:readdata -> mm_interconnect_0:altpll_mipi_pll_slave_readdata
	wire    [1:0] mm_interconnect_0_altpll_mipi_pll_slave_address;           // mm_interconnect_0:altpll_mipi_pll_slave_address -> altpll_mipi:address
	wire          mm_interconnect_0_altpll_mipi_pll_slave_read;              // mm_interconnect_0:altpll_mipi_pll_slave_read -> altpll_mipi:read
	wire          mm_interconnect_0_altpll_mipi_pll_slave_write;             // mm_interconnect_0:altpll_mipi_pll_slave_write -> altpll_mipi:write
	wire   [31:0] mm_interconnect_0_altpll_mipi_pll_slave_writedata;         // mm_interconnect_0:altpll_mipi_pll_slave_writedata -> altpll_mipi:writedata
	wire          mm_interconnect_0_timer_s1_chipselect;                     // mm_interconnect_0:timer_s1_chipselect -> timer:chipselect
	wire   [15:0] mm_interconnect_0_timer_s1_readdata;                       // timer:readdata -> mm_interconnect_0:timer_s1_readdata
	wire    [2:0] mm_interconnect_0_timer_s1_address;                        // mm_interconnect_0:timer_s1_address -> timer:address
	wire          mm_interconnect_0_timer_s1_write;                          // mm_interconnect_0:timer_s1_write -> timer:write_n
	wire   [15:0] mm_interconnect_0_timer_s1_writedata;                      // mm_interconnect_0:timer_s1_writedata -> timer:writedata
	wire          mm_interconnect_0_led_s1_chipselect;                       // mm_interconnect_0:led_s1_chipselect -> led:chipselect
	wire   [31:0] mm_interconnect_0_led_s1_readdata;                         // led:readdata -> mm_interconnect_0:led_s1_readdata
	wire    [1:0] mm_interconnect_0_led_s1_address;                          // mm_interconnect_0:led_s1_address -> led:address
	wire          mm_interconnect_0_led_s1_write;                            // mm_interconnect_0:led_s1_write -> led:write_n
	wire   [31:0] mm_interconnect_0_led_s1_writedata;                        // mm_interconnect_0:led_s1_writedata -> led:writedata
	wire   [31:0] mm_interconnect_0_sw_s1_readdata;                          // sw:readdata -> mm_interconnect_0:sw_s1_readdata
	wire    [1:0] mm_interconnect_0_sw_s1_address;                           // mm_interconnect_0:sw_s1_address -> sw:address
	wire   [31:0] mm_interconnect_0_ddr3_status_s1_readdata;                 // ddr3_status:readdata -> mm_interconnect_0:ddr3_status_s1_readdata
	wire    [1:0] mm_interconnect_0_ddr3_status_s1_address;                  // mm_interconnect_0:ddr3_status_s1_address -> ddr3_status:address
	wire          irq_mapper_receiver1_irq;                                  // jtag_uart:av_irq -> irq_mapper:receiver1_irq
	wire          irq_mapper_receiver2_irq;                                  // timer:irq -> irq_mapper:receiver2_irq
	wire   [31:0] nios2_gen2_irq_irq;                                        // irq_mapper:sender_irq -> nios2_gen2:irq
	wire          irq_mapper_receiver0_irq;                                  // irq_synchronizer:sender_irq -> irq_mapper:receiver0_irq
	wire    [0:0] irq_synchronizer_receiver_irq;                             // alt_vip_vfr_1:slave_irq -> irq_synchronizer:receiver_irq
	wire          irq_mapper_receiver3_irq;                                  // irq_synchronizer_001:sender_irq -> irq_mapper:receiver3_irq
	wire    [0:0] irq_synchronizer_001_receiver_irq;                         // hdmi_cvo:status_update_irq_irq -> irq_synchronizer_001:receiver_irq
	wire          rst_controller_reset_out_reset;                            // rst_controller:reset_out -> [alt_vip_cpr_1:reset, alt_vip_vfr_1:reset, irq_synchronizer:receiver_reset, mm_interconnect_0:alt_vip_vfr_1_clock_reset_reset_reset_bridge_in_reset_reset]
	wire          rst_controller_001_reset_out_reset;                        // rst_controller_001:reset_out -> [alt_vip_vfr_1:master_reset, mm_interconnect_0:alt_vip_vfr_1_clock_master_reset_reset_bridge_in_reset_reset]
	wire          rst_controller_002_reset_out_reset;                        // rst_controller_002:reset_out -> [altpll_mipi:reset, altpll_sys:reset, mm_interconnect_0:altpll_mipi_inclk_interface_reset_reset_bridge_in_reset_reset]
	wire          rst_controller_003_reset_out_reset;                        // rst_controller_003:reset_out -> [hdmi_cvo:main_reset_reset, irq_synchronizer_001:receiver_reset]
	wire          rst_controller_004_reset_out_reset;                        // rst_controller_004:reset_out -> [jtag_uart:rst_n, mm_interconnect_0:onchip_memory2_reset1_reset_bridge_in_reset_reset, onchip_memory2:reset, rst_translator:in_reset, sysid_qsys:reset_n, timer:reset_n]
	wire          rst_controller_004_reset_out_reset_req;                    // rst_controller_004:reset_req -> [onchip_memory2:reset_req, rst_translator:reset_req_in]
	wire          rst_controller_005_reset_out_reset;                        // rst_controller_005:reset_out -> [led:reset_n, mm_interconnect_0:led_reset_reset_bridge_in_reset_reset, sw:reset_n]
	wire          rst_controller_006_reset_out_reset;                        // rst_controller_006:reset_out -> [irq_mapper:reset, irq_synchronizer:sender_reset, irq_synchronizer_001:sender_reset, mm_interconnect_0:nios2_gen2_reset_reset_bridge_in_reset_reset, nios2_gen2:reset_n, rst_translator_001:in_reset]
	wire          rst_controller_006_reset_out_reset_req;                    // rst_controller_006:reset_req -> [nios2_gen2:reset_req, rst_translator_001:reset_req_in]
	wire          rst_controller_007_reset_out_reset;                        // rst_controller_007:reset_out -> [mm_interconnect_0:mem_if_ddr3_emif_avl_translator_reset_reset_bridge_in_reset_reset, mm_interconnect_0:mem_if_ddr3_emif_soft_reset_reset_bridge_in_reset_reset]

	deca_vip_alt_vip_cpr_1 alt_vip_cpr_1 (
		.clock               (altpll_sys_c1_clk),                                   // clock.clk
		.reset               (rst_controller_reset_out_reset),                      // reset.reset
		.din0_ready          (alt_vip_vfr_1_avalon_streaming_source_ready),         //  din0.ready
		.din0_valid          (alt_vip_vfr_1_avalon_streaming_source_valid),         //      .valid
		.din0_data           (alt_vip_vfr_1_avalon_streaming_source_data),          //      .data
		.din0_startofpacket  (alt_vip_vfr_1_avalon_streaming_source_startofpacket), //      .startofpacket
		.din0_endofpacket    (alt_vip_vfr_1_avalon_streaming_source_endofpacket),   //      .endofpacket
		.dout0_ready         (alt_vip_cpr_1_dout0_ready),                           // dout0.ready
		.dout0_valid         (alt_vip_cpr_1_dout0_valid),                           //      .valid
		.dout0_data          (alt_vip_cpr_1_dout0_data),                            //      .data
		.dout0_startofpacket (alt_vip_cpr_1_dout0_startofpacket),                   //      .startofpacket
		.dout0_endofpacket   (alt_vip_cpr_1_dout0_endofpacket)                      //      .endofpacket
	);

	alt_vipvfr131_vfr #(
		.BITS_PER_PIXEL_PER_COLOR_PLANE (8),
		.NUMBER_OF_CHANNELS_IN_PARALLEL (4),
		.NUMBER_OF_CHANNELS_IN_SEQUENCE (1),
		.MAX_IMAGE_WIDTH                (1280),
		.MAX_IMAGE_HEIGHT               (800),
		.MEM_PORT_WIDTH                 (256),
		.RMASTER_FIFO_DEPTH             (1024),
		.RMASTER_BURST_TARGET           (32),
		.CLOCKS_ARE_SEPARATE            (1)
	) alt_vip_vfr_1 (
		.clock                (altpll_sys_c1_clk),                                      //             clock_reset.clk
		.reset                (rst_controller_reset_out_reset),                         //       clock_reset_reset.reset
		.master_clock         (altpll_sys_c1_clk),                                      //            clock_master.clk
		.master_reset         (rst_controller_001_reset_out_reset),                     //      clock_master_reset.reset
		.slave_address        (mm_interconnect_0_alt_vip_vfr_1_avalon_slave_address),   //            avalon_slave.address
		.slave_write          (mm_interconnect_0_alt_vip_vfr_1_avalon_slave_write),     //                        .write
		.slave_writedata      (mm_interconnect_0_alt_vip_vfr_1_avalon_slave_writedata), //                        .writedata
		.slave_read           (mm_interconnect_0_alt_vip_vfr_1_avalon_slave_read),      //                        .read
		.slave_readdata       (mm_interconnect_0_alt_vip_vfr_1_avalon_slave_readdata),  //                        .readdata
		.slave_irq            (irq_synchronizer_receiver_irq),                          //        interrupt_sender.irq
		.dout_data            (alt_vip_vfr_1_avalon_streaming_source_data),             // avalon_streaming_source.data
		.dout_valid           (alt_vip_vfr_1_avalon_streaming_source_valid),            //                        .valid
		.dout_ready           (alt_vip_vfr_1_avalon_streaming_source_ready),            //                        .ready
		.dout_startofpacket   (alt_vip_vfr_1_avalon_streaming_source_startofpacket),    //                        .startofpacket
		.dout_endofpacket     (alt_vip_vfr_1_avalon_streaming_source_endofpacket),      //                        .endofpacket
		.master_address       (alt_vip_vfr_1_avalon_master_address),                    //           avalon_master.address
		.master_burstcount    (alt_vip_vfr_1_avalon_master_burstcount),                 //                        .burstcount
		.master_readdata      (alt_vip_vfr_1_avalon_master_readdata),                   //                        .readdata
		.master_read          (alt_vip_vfr_1_avalon_master_read),                       //                        .read
		.master_readdatavalid (alt_vip_vfr_1_avalon_master_readdatavalid),              //                        .readdatavalid
		.master_waitrequest   (alt_vip_vfr_1_avalon_master_waitrequest)                 //                        .waitrequest
	);

	deca_vip_altpll_mipi altpll_mipi (
		.clk       (clk_clk),                                           //       inclk_interface.clk
		.reset     (rst_controller_002_reset_out_reset),                // inclk_interface_reset.reset
		.read      (mm_interconnect_0_altpll_mipi_pll_slave_read),      //             pll_slave.read
		.write     (mm_interconnect_0_altpll_mipi_pll_slave_write),     //                      .write
		.address   (mm_interconnect_0_altpll_mipi_pll_slave_address),   //                      .address
		.readdata  (mm_interconnect_0_altpll_mipi_pll_slave_readdata),  //                      .readdata
		.writedata (mm_interconnect_0_altpll_mipi_pll_slave_writedata), //                      .writedata
		.c0        (altpll_mipi_clk_clk),                               //                    c0.clk
		.areset    (),                                                  //        areset_conduit.export
		.locked    (),                                                  //        locked_conduit.export
		.phasedone ()                                                   //     phasedone_conduit.export
	);

	deca_vip_altpll_sys altpll_sys (
		.clk       (clk_clk),                            //       inclk_interface.clk
		.reset     (rst_controller_002_reset_out_reset), // inclk_interface_reset.reset
		.read      (),                                   //             pll_slave.read
		.write     (),                                   //                      .write
		.address   (),                                   //                      .address
		.readdata  (),                                   //                      .readdata
		.writedata (),                                   //                      .writedata
		.c0        (clock_bridge_vip_out_clk_clk),       //                    c0.clk
		.c1        (altpll_sys_c1_clk),                  //                    c1.clk
		.c2        (altpll_sys_hdmi_clk),                //                    c2.clk
		.areset    (),                                   //        areset_conduit.export
		.locked    (),                                   //        locked_conduit.export
		.phasedone ()                                    //     phasedone_conduit.export
	);

	deca_vip_ddr3_status ddr3_status (
		.clk      (clock_bridge_vip_out_clk_clk),              //                 clk.clk
		.reset_n  (~nios2_gen2_debug_reset_request_reset),     //               reset.reset_n
		.address  (mm_interconnect_0_ddr3_status_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_ddr3_status_s1_readdata), //                    .readdata
		.in_port  (ddr3_status_external_connection_export)     // external_connection.export
	);

	deca_vip_hdmi_cvo #(
		.NUMBER_OF_COLOUR_PLANES       (3),
		.COLOUR_PLANES_ARE_IN_PARALLEL (1),
		.BPS                           (8),
		.INTERLACED                    (0),
		.H_ACTIVE_PIXELS               (1280),
		.V_ACTIVE_LINES                (800),
		.ACCEPT_COLOURS_IN_SEQ         (0),
		.FIFO_DEPTH                    (1280),
		.CLOCKS_ARE_SAME               (0),
		.USE_CONTROL                   (0),
		.NO_OF_MODES                   (1),
		.THRESHOLD                     (1279),
		.STD_WIDTH                     (1),
		.GENERATE_SYNC                 (0),
		.USE_EMBEDDED_SYNCS            (0),
		.AP_LINE                       (0),
		.V_BLANK                       (0),
		.H_BLANK                       (0),
		.H_SYNC_LENGTH                 (136),
		.H_FRONT_PORCH                 (64),
		.H_BACK_PORCH                  (200),
		.V_SYNC_LENGTH                 (3),
		.V_FRONT_PORCH                 (1),
		.V_BACK_PORCH                  (24),
		.F_RISING_EDGE                 (0),
		.F_FALLING_EDGE                (0),
		.FIELD0_V_RISING_EDGE          (0),
		.FIELD0_V_BLANK                (0),
		.FIELD0_V_SYNC_LENGTH          (0),
		.FIELD0_V_FRONT_PORCH          (0),
		.FIELD0_V_BACK_PORCH           (0),
		.ANC_LINE                      (0),
		.FIELD0_ANC_LINE               (0),
		.SRC_WIDTH                     (8),
		.DST_WIDTH                     (8),
		.CONTEXT_WIDTH                 (8),
		.TASK_WIDTH                    (8)
	) hdmi_cvo (
		.clocked_video_vid_clk       (hdmi_cvo_vid_clk),                   //     clocked_video.vid_clk
		.clocked_video_vid_data      (hdmi_cvo_vid_data),                  //                  .vid_data
		.clocked_video_underflow     (hdmi_cvo_underflow),                 //                  .underflow
		.clocked_video_vid_datavalid (hdmi_cvo_vid_datavalid),             //                  .vid_datavalid
		.clocked_video_vid_v_sync    (hdmi_cvo_vid_v_sync),                //                  .vid_v_sync
		.clocked_video_vid_h_sync    (hdmi_cvo_vid_h_sync),                //                  .vid_h_sync
		.clocked_video_vid_f         (hdmi_cvo_vid_f),                     //                  .vid_f
		.clocked_video_vid_h         (hdmi_cvo_vid_h),                     //                  .vid_h
		.clocked_video_vid_v         (hdmi_cvo_vid_v),                     //                  .vid_v
		.main_clock_clk              (altpll_sys_c1_clk),                  //        main_clock.clk
		.main_reset_reset            (rst_controller_003_reset_out_reset), //        main_reset.reset
		.din_data                    (alt_vip_cpr_1_dout0_data),           //               din.data
		.din_valid                   (alt_vip_cpr_1_dout0_valid),          //                  .valid
		.din_startofpacket           (alt_vip_cpr_1_dout0_startofpacket),  //                  .startofpacket
		.din_endofpacket             (alt_vip_cpr_1_dout0_endofpacket),    //                  .endofpacket
		.din_ready                   (alt_vip_cpr_1_dout0_ready),          //                  .ready
		.status_update_irq_irq       (irq_synchronizer_001_receiver_irq)   // status_update_irq.irq
	);

	deca_vip_jtag_uart jtag_uart (
		.clk            (clock_bridge_vip_out_clk_clk),                              //               clk.clk
		.rst_n          (~rst_controller_004_reset_out_reset),                       //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver1_irq)                                   //               irq.irq
	);

	deca_vip_led led (
		.clk        (clk_clk),                             //                 clk.clk
		.reset_n    (~rst_controller_005_reset_out_reset), //               reset.reset_n
		.address    (mm_interconnect_0_led_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_led_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_led_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_led_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_led_s1_readdata),   //                    .readdata
		.out_port   (led_external_connection_export)       // external_connection.export
	);

	deca_vip_mem_if_ddr3_emif mem_if_ddr3_emif (
		.pll_ref_clk        (mem_if_ddr3_emif_pll_ref_clk_clk),                          //      pll_ref_clk.clk
		.global_reset_n     (~nios2_gen2_debug_reset_request_reset),                     //     global_reset.reset_n
		.soft_reset_n       (~nios2_gen2_debug_reset_request_reset),                     //       soft_reset.reset_n
		.afi_clk            (mem_if_ddr3_emif_afi_clk_clk),                              //          afi_clk.clk
		.afi_half_clk       (),                                                          //     afi_half_clk.clk
		.afi_reset_n        (),                                                          //        afi_reset.reset_n
		.afi_reset_export_n (),                                                          // afi_reset_export.reset_n
		.mem_a              (memory_mem_a),                                              //           memory.mem_a
		.mem_ba             (memory_mem_ba),                                             //                 .mem_ba
		.mem_ck             (memory_mem_ck),                                             //                 .mem_ck
		.mem_ck_n           (memory_mem_ck_n),                                           //                 .mem_ck_n
		.mem_cke            (memory_mem_cke),                                            //                 .mem_cke
		.mem_cs_n           (memory_mem_cs_n),                                           //                 .mem_cs_n
		.mem_dm             (memory_mem_dm),                                             //                 .mem_dm
		.mem_ras_n          (memory_mem_ras_n),                                          //                 .mem_ras_n
		.mem_cas_n          (memory_mem_cas_n),                                          //                 .mem_cas_n
		.mem_we_n           (memory_mem_we_n),                                           //                 .mem_we_n
		.mem_reset_n        (memory_mem_reset_n),                                        //                 .mem_reset_n
		.mem_dq             (memory_mem_dq),                                             //                 .mem_dq
		.mem_dqs            (memory_mem_dqs),                                            //                 .mem_dqs
		.mem_dqs_n          (memory_mem_dqs_n),                                          //                 .mem_dqs_n
		.mem_odt            (memory_mem_odt),                                            //                 .mem_odt
		.avl_ready          (mm_interconnect_0_mem_if_ddr3_emif_avl_waitrequest),        //              avl.waitrequest_n
		.avl_burstbegin     (mm_interconnect_0_mem_if_ddr3_emif_avl_beginbursttransfer), //                 .beginbursttransfer
		.avl_addr           (mm_interconnect_0_mem_if_ddr3_emif_avl_address),            //                 .address
		.avl_rdata_valid    (mm_interconnect_0_mem_if_ddr3_emif_avl_readdatavalid),      //                 .readdatavalid
		.avl_rdata          (mm_interconnect_0_mem_if_ddr3_emif_avl_readdata),           //                 .readdata
		.avl_wdata          (mm_interconnect_0_mem_if_ddr3_emif_avl_writedata),          //                 .writedata
		.avl_be             (mm_interconnect_0_mem_if_ddr3_emif_avl_byteenable),         //                 .byteenable
		.avl_read_req       (mm_interconnect_0_mem_if_ddr3_emif_avl_read),               //                 .read
		.avl_write_req      (mm_interconnect_0_mem_if_ddr3_emif_avl_write),              //                 .write
		.avl_size           (mm_interconnect_0_mem_if_ddr3_emif_avl_burstcount),         //                 .burstcount
		.local_init_done    (mem_if_ddr3_emif_status_local_init_done),                   //           status.local_init_done
		.local_cal_success  (mem_if_ddr3_emif_status_local_cal_success),                 //                 .local_cal_success
		.local_cal_fail     (mem_if_ddr3_emif_status_local_cal_fail),                    //                 .local_cal_fail
		.pll_mem_clk        (mem_if_ddr3_emif_pll_sharing_pll_mem_clk),                  //      pll_sharing.pll_mem_clk
		.pll_write_clk      (mem_if_ddr3_emif_pll_sharing_pll_write_clk),                //                 .pll_write_clk
		.pll_locked         (mem_if_ddr3_emif_pll_sharing_pll_locked),                   //                 .pll_locked
		.pll_capture0_clk   (mem_if_ddr3_emif_pll_sharing_pll_capture0_clk),             //                 .pll_capture0_clk
		.pll_capture1_clk   (mem_if_ddr3_emif_pll_sharing_pll_capture1_clk)              //                 .pll_capture1_clk
	);

	deca_vip_nios2_gen2 nios2_gen2 (
		.clk                                 (clock_bridge_vip_out_clk_clk),                             //                       clk.clk
		.reset_n                             (~rst_controller_006_reset_out_reset),                      //                     reset.reset_n
		.reset_req                           (rst_controller_006_reset_out_reset_req),                   //                          .reset_req
		.d_address                           (nios2_gen2_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios2_gen2_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios2_gen2_data_master_read),                              //                          .read
		.d_readdata                          (nios2_gen2_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios2_gen2_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios2_gen2_data_master_write),                             //                          .write
		.d_writedata                         (nios2_gen2_data_master_writedata),                         //                          .writedata
		.d_readdatavalid                     (nios2_gen2_data_master_readdatavalid),                     //                          .readdatavalid
		.debug_mem_slave_debugaccess_to_roms (nios2_gen2_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios2_gen2_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios2_gen2_instruction_master_read),                       //                          .read
		.i_readdata                          (nios2_gen2_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios2_gen2_instruction_master_waitrequest),                //                          .waitrequest
		.i_readdatavalid                     (nios2_gen2_instruction_master_readdatavalid),              //                          .readdatavalid
		.irq                                 (nios2_gen2_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (nios2_gen2_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios2_gen2_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios2_gen2_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios2_gen2_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios2_gen2_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios2_gen2_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios2_gen2_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios2_gen2_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios2_gen2_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                          // custom_instruction_master.readra
	);

	deca_vip_onchip_memory2 onchip_memory2 (
		.clk        (clock_bridge_vip_out_clk_clk),                   //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory2_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory2_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory2_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory2_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory2_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory2_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory2_s1_byteenable), //       .byteenable
		.reset      (rst_controller_004_reset_out_reset),             // reset1.reset
		.reset_req  (rst_controller_004_reset_out_reset_req)          //       .reset_req
	);

	deca_vip_sw sw (
		.clk      (clk_clk),                             //                 clk.clk
		.reset_n  (~rst_controller_005_reset_out_reset), //               reset.reset_n
		.address  (mm_interconnect_0_sw_s1_address),     //                  s1.address
		.readdata (mm_interconnect_0_sw_s1_readdata),    //                    .readdata
		.in_port  (sw_external_connection_export)        // external_connection.export
	);

	deca_vip_sysid_qsys sysid_qsys (
		.clock    (clock_bridge_vip_out_clk_clk),                        //           clk.clk
		.reset_n  (~rst_controller_004_reset_out_reset),                 //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_qsys_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_qsys_control_slave_address)   //              .address
	);

	deca_vip_timer timer (
		.clk        (clock_bridge_vip_out_clk_clk),          //   clk.clk
		.reset_n    (~rst_controller_004_reset_out_reset),   // reset.reset_n
		.address    (mm_interconnect_0_timer_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver2_irq)               //   irq.irq
	);

	deca_vip_mm_interconnect_0 mm_interconnect_0 (
		.altpll_sys_c0_clk                                                 (clock_bridge_vip_out_clk_clk),                              //                                               altpll_sys_c0.clk
		.altpll_sys_c1_clk                                                 (altpll_sys_c1_clk),                                         //                                               altpll_sys_c1.clk
		.clk_50_clk_clk                                                    (clk_clk),                                                   //                                                  clk_50_clk.clk
		.mem_if_ddr3_emif_afi_clk_clk                                      (mem_if_ddr3_emif_afi_clk_clk),                              //                                    mem_if_ddr3_emif_afi_clk.clk
		.alt_vip_vfr_1_clock_master_reset_reset_bridge_in_reset_reset      (rst_controller_001_reset_out_reset),                        //      alt_vip_vfr_1_clock_master_reset_reset_bridge_in_reset.reset
		.alt_vip_vfr_1_clock_reset_reset_reset_bridge_in_reset_reset       (rst_controller_reset_out_reset),                            //       alt_vip_vfr_1_clock_reset_reset_reset_bridge_in_reset.reset
		.altpll_mipi_inclk_interface_reset_reset_bridge_in_reset_reset     (rst_controller_002_reset_out_reset),                        //     altpll_mipi_inclk_interface_reset_reset_bridge_in_reset.reset
		.ddr3_status_reset_reset_bridge_in_reset_reset                     (nios2_gen2_debug_reset_request_reset),                      //                     ddr3_status_reset_reset_bridge_in_reset.reset
		.led_reset_reset_bridge_in_reset_reset                             (rst_controller_005_reset_out_reset),                        //                             led_reset_reset_bridge_in_reset.reset
		.mem_if_ddr3_emif_avl_translator_reset_reset_bridge_in_reset_reset (rst_controller_007_reset_out_reset),                        // mem_if_ddr3_emif_avl_translator_reset_reset_bridge_in_reset.reset
		.mem_if_ddr3_emif_soft_reset_reset_bridge_in_reset_reset           (rst_controller_007_reset_out_reset),                        //           mem_if_ddr3_emif_soft_reset_reset_bridge_in_reset.reset
		.nios2_gen2_reset_reset_bridge_in_reset_reset                      (rst_controller_006_reset_out_reset),                        //                      nios2_gen2_reset_reset_bridge_in_reset.reset
		.onchip_memory2_reset1_reset_bridge_in_reset_reset                 (rst_controller_004_reset_out_reset),                        //                 onchip_memory2_reset1_reset_bridge_in_reset.reset
		.alt_vip_vfr_1_avalon_master_address                               (alt_vip_vfr_1_avalon_master_address),                       //                                 alt_vip_vfr_1_avalon_master.address
		.alt_vip_vfr_1_avalon_master_waitrequest                           (alt_vip_vfr_1_avalon_master_waitrequest),                   //                                                            .waitrequest
		.alt_vip_vfr_1_avalon_master_burstcount                            (alt_vip_vfr_1_avalon_master_burstcount),                    //                                                            .burstcount
		.alt_vip_vfr_1_avalon_master_read                                  (alt_vip_vfr_1_avalon_master_read),                          //                                                            .read
		.alt_vip_vfr_1_avalon_master_readdata                              (alt_vip_vfr_1_avalon_master_readdata),                      //                                                            .readdata
		.alt_vip_vfr_1_avalon_master_readdatavalid                         (alt_vip_vfr_1_avalon_master_readdatavalid),                 //                                                            .readdatavalid
		.nios2_gen2_data_master_address                                    (nios2_gen2_data_master_address),                            //                                      nios2_gen2_data_master.address
		.nios2_gen2_data_master_waitrequest                                (nios2_gen2_data_master_waitrequest),                        //                                                            .waitrequest
		.nios2_gen2_data_master_byteenable                                 (nios2_gen2_data_master_byteenable),                         //                                                            .byteenable
		.nios2_gen2_data_master_read                                       (nios2_gen2_data_master_read),                               //                                                            .read
		.nios2_gen2_data_master_readdata                                   (nios2_gen2_data_master_readdata),                           //                                                            .readdata
		.nios2_gen2_data_master_readdatavalid                              (nios2_gen2_data_master_readdatavalid),                      //                                                            .readdatavalid
		.nios2_gen2_data_master_write                                      (nios2_gen2_data_master_write),                              //                                                            .write
		.nios2_gen2_data_master_writedata                                  (nios2_gen2_data_master_writedata),                          //                                                            .writedata
		.nios2_gen2_data_master_debugaccess                                (nios2_gen2_data_master_debugaccess),                        //                                                            .debugaccess
		.nios2_gen2_instruction_master_address                             (nios2_gen2_instruction_master_address),                     //                               nios2_gen2_instruction_master.address
		.nios2_gen2_instruction_master_waitrequest                         (nios2_gen2_instruction_master_waitrequest),                 //                                                            .waitrequest
		.nios2_gen2_instruction_master_read                                (nios2_gen2_instruction_master_read),                        //                                                            .read
		.nios2_gen2_instruction_master_readdata                            (nios2_gen2_instruction_master_readdata),                    //                                                            .readdata
		.nios2_gen2_instruction_master_readdatavalid                       (nios2_gen2_instruction_master_readdatavalid),               //                                                            .readdatavalid
		.alt_vip_vfr_1_avalon_slave_address                                (mm_interconnect_0_alt_vip_vfr_1_avalon_slave_address),      //                                  alt_vip_vfr_1_avalon_slave.address
		.alt_vip_vfr_1_avalon_slave_write                                  (mm_interconnect_0_alt_vip_vfr_1_avalon_slave_write),        //                                                            .write
		.alt_vip_vfr_1_avalon_slave_read                                   (mm_interconnect_0_alt_vip_vfr_1_avalon_slave_read),         //                                                            .read
		.alt_vip_vfr_1_avalon_slave_readdata                               (mm_interconnect_0_alt_vip_vfr_1_avalon_slave_readdata),     //                                                            .readdata
		.alt_vip_vfr_1_avalon_slave_writedata                              (mm_interconnect_0_alt_vip_vfr_1_avalon_slave_writedata),    //                                                            .writedata
		.altpll_mipi_pll_slave_address                                     (mm_interconnect_0_altpll_mipi_pll_slave_address),           //                                       altpll_mipi_pll_slave.address
		.altpll_mipi_pll_slave_write                                       (mm_interconnect_0_altpll_mipi_pll_slave_write),             //                                                            .write
		.altpll_mipi_pll_slave_read                                        (mm_interconnect_0_altpll_mipi_pll_slave_read),              //                                                            .read
		.altpll_mipi_pll_slave_readdata                                    (mm_interconnect_0_altpll_mipi_pll_slave_readdata),          //                                                            .readdata
		.altpll_mipi_pll_slave_writedata                                   (mm_interconnect_0_altpll_mipi_pll_slave_writedata),         //                                                            .writedata
		.ddr3_status_s1_address                                            (mm_interconnect_0_ddr3_status_s1_address),                  //                                              ddr3_status_s1.address
		.ddr3_status_s1_readdata                                           (mm_interconnect_0_ddr3_status_s1_readdata),                 //                                                            .readdata
		.jtag_uart_avalon_jtag_slave_address                               (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                                 jtag_uart_avalon_jtag_slave.address
		.jtag_uart_avalon_jtag_slave_write                                 (mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),       //                                                            .write
		.jtag_uart_avalon_jtag_slave_read                                  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),        //                                                            .read
		.jtag_uart_avalon_jtag_slave_readdata                              (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                                                            .readdata
		.jtag_uart_avalon_jtag_slave_writedata                             (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                                                            .writedata
		.jtag_uart_avalon_jtag_slave_waitrequest                           (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                                                            .waitrequest
		.jtag_uart_avalon_jtag_slave_chipselect                            (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  //                                                            .chipselect
		.led_s1_address                                                    (mm_interconnect_0_led_s1_address),                          //                                                      led_s1.address
		.led_s1_write                                                      (mm_interconnect_0_led_s1_write),                            //                                                            .write
		.led_s1_readdata                                                   (mm_interconnect_0_led_s1_readdata),                         //                                                            .readdata
		.led_s1_writedata                                                  (mm_interconnect_0_led_s1_writedata),                        //                                                            .writedata
		.led_s1_chipselect                                                 (mm_interconnect_0_led_s1_chipselect),                       //                                                            .chipselect
		.mem_if_ddr3_emif_avl_address                                      (mm_interconnect_0_mem_if_ddr3_emif_avl_address),            //                                        mem_if_ddr3_emif_avl.address
		.mem_if_ddr3_emif_avl_write                                        (mm_interconnect_0_mem_if_ddr3_emif_avl_write),              //                                                            .write
		.mem_if_ddr3_emif_avl_read                                         (mm_interconnect_0_mem_if_ddr3_emif_avl_read),               //                                                            .read
		.mem_if_ddr3_emif_avl_readdata                                     (mm_interconnect_0_mem_if_ddr3_emif_avl_readdata),           //                                                            .readdata
		.mem_if_ddr3_emif_avl_writedata                                    (mm_interconnect_0_mem_if_ddr3_emif_avl_writedata),          //                                                            .writedata
		.mem_if_ddr3_emif_avl_beginbursttransfer                           (mm_interconnect_0_mem_if_ddr3_emif_avl_beginbursttransfer), //                                                            .beginbursttransfer
		.mem_if_ddr3_emif_avl_burstcount                                   (mm_interconnect_0_mem_if_ddr3_emif_avl_burstcount),         //                                                            .burstcount
		.mem_if_ddr3_emif_avl_byteenable                                   (mm_interconnect_0_mem_if_ddr3_emif_avl_byteenable),         //                                                            .byteenable
		.mem_if_ddr3_emif_avl_readdatavalid                                (mm_interconnect_0_mem_if_ddr3_emif_avl_readdatavalid),      //                                                            .readdatavalid
		.mem_if_ddr3_emif_avl_waitrequest                                  (~mm_interconnect_0_mem_if_ddr3_emif_avl_waitrequest),       //                                                            .waitrequest
		.nios2_gen2_debug_mem_slave_address                                (mm_interconnect_0_nios2_gen2_debug_mem_slave_address),      //                                  nios2_gen2_debug_mem_slave.address
		.nios2_gen2_debug_mem_slave_write                                  (mm_interconnect_0_nios2_gen2_debug_mem_slave_write),        //                                                            .write
		.nios2_gen2_debug_mem_slave_read                                   (mm_interconnect_0_nios2_gen2_debug_mem_slave_read),         //                                                            .read
		.nios2_gen2_debug_mem_slave_readdata                               (mm_interconnect_0_nios2_gen2_debug_mem_slave_readdata),     //                                                            .readdata
		.nios2_gen2_debug_mem_slave_writedata                              (mm_interconnect_0_nios2_gen2_debug_mem_slave_writedata),    //                                                            .writedata
		.nios2_gen2_debug_mem_slave_byteenable                             (mm_interconnect_0_nios2_gen2_debug_mem_slave_byteenable),   //                                                            .byteenable
		.nios2_gen2_debug_mem_slave_waitrequest                            (mm_interconnect_0_nios2_gen2_debug_mem_slave_waitrequest),  //                                                            .waitrequest
		.nios2_gen2_debug_mem_slave_debugaccess                            (mm_interconnect_0_nios2_gen2_debug_mem_slave_debugaccess),  //                                                            .debugaccess
		.onchip_memory2_s1_address                                         (mm_interconnect_0_onchip_memory2_s1_address),               //                                           onchip_memory2_s1.address
		.onchip_memory2_s1_write                                           (mm_interconnect_0_onchip_memory2_s1_write),                 //                                                            .write
		.onchip_memory2_s1_readdata                                        (mm_interconnect_0_onchip_memory2_s1_readdata),              //                                                            .readdata
		.onchip_memory2_s1_writedata                                       (mm_interconnect_0_onchip_memory2_s1_writedata),             //                                                            .writedata
		.onchip_memory2_s1_byteenable                                      (mm_interconnect_0_onchip_memory2_s1_byteenable),            //                                                            .byteenable
		.onchip_memory2_s1_chipselect                                      (mm_interconnect_0_onchip_memory2_s1_chipselect),            //                                                            .chipselect
		.onchip_memory2_s1_clken                                           (mm_interconnect_0_onchip_memory2_s1_clken),                 //                                                            .clken
		.sw_s1_address                                                     (mm_interconnect_0_sw_s1_address),                           //                                                       sw_s1.address
		.sw_s1_readdata                                                    (mm_interconnect_0_sw_s1_readdata),                          //                                                            .readdata
		.sysid_qsys_control_slave_address                                  (mm_interconnect_0_sysid_qsys_control_slave_address),        //                                    sysid_qsys_control_slave.address
		.sysid_qsys_control_slave_readdata                                 (mm_interconnect_0_sysid_qsys_control_slave_readdata),       //                                                            .readdata
		.timer_s1_address                                                  (mm_interconnect_0_timer_s1_address),                        //                                                    timer_s1.address
		.timer_s1_write                                                    (mm_interconnect_0_timer_s1_write),                          //                                                            .write
		.timer_s1_readdata                                                 (mm_interconnect_0_timer_s1_readdata),                       //                                                            .readdata
		.timer_s1_writedata                                                (mm_interconnect_0_timer_s1_writedata),                      //                                                            .writedata
		.timer_s1_chipselect                                               (mm_interconnect_0_timer_s1_chipselect)                      //                                                            .chipselect
	);

	deca_vip_irq_mapper irq_mapper (
		.clk           (clock_bridge_vip_out_clk_clk),       //       clk.clk
		.reset         (rst_controller_006_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),           // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),           // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),           // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),           // receiver3.irq
		.sender_irq    (nios2_gen2_irq_irq)                  //    sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer (
		.receiver_clk   (altpll_sys_c1_clk),                  //       receiver_clk.clk
		.sender_clk     (clock_bridge_vip_out_clk_clk),       //         sender_clk.clk
		.receiver_reset (rst_controller_reset_out_reset),     // receiver_clk_reset.reset
		.sender_reset   (rst_controller_006_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_receiver_irq),      //           receiver.irq
		.sender_irq     (irq_mapper_receiver0_irq)            //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_001 (
		.receiver_clk   (altpll_sys_c1_clk),                  //       receiver_clk.clk
		.sender_clk     (clock_bridge_vip_out_clk_clk),       //         sender_clk.clk
		.receiver_reset (rst_controller_003_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_006_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_001_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver3_irq)            //             sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (nios2_gen2_debug_reset_request_reset), // reset_in0.reset
		.clk            (altpll_sys_c1_clk),                    //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),       // reset_out.reset
		.reset_req      (),                                     // (terminated)
		.reset_req_in0  (1'b0),                                 // (terminated)
		.reset_in1      (1'b0),                                 // (terminated)
		.reset_req_in1  (1'b0),                                 // (terminated)
		.reset_in2      (1'b0),                                 // (terminated)
		.reset_req_in2  (1'b0),                                 // (terminated)
		.reset_in3      (1'b0),                                 // (terminated)
		.reset_req_in3  (1'b0),                                 // (terminated)
		.reset_in4      (1'b0),                                 // (terminated)
		.reset_req_in4  (1'b0),                                 // (terminated)
		.reset_in5      (1'b0),                                 // (terminated)
		.reset_req_in5  (1'b0),                                 // (terminated)
		.reset_in6      (1'b0),                                 // (terminated)
		.reset_req_in6  (1'b0),                                 // (terminated)
		.reset_in7      (1'b0),                                 // (terminated)
		.reset_req_in7  (1'b0),                                 // (terminated)
		.reset_in8      (1'b0),                                 // (terminated)
		.reset_req_in8  (1'b0),                                 // (terminated)
		.reset_in9      (1'b0),                                 // (terminated)
		.reset_req_in9  (1'b0),                                 // (terminated)
		.reset_in10     (1'b0),                                 // (terminated)
		.reset_req_in10 (1'b0),                                 // (terminated)
		.reset_in11     (1'b0),                                 // (terminated)
		.reset_req_in11 (1'b0),                                 // (terminated)
		.reset_in12     (1'b0),                                 // (terminated)
		.reset_req_in12 (1'b0),                                 // (terminated)
		.reset_in13     (1'b0),                                 // (terminated)
		.reset_req_in13 (1'b0),                                 // (terminated)
		.reset_in14     (1'b0),                                 // (terminated)
		.reset_req_in14 (1'b0),                                 // (terminated)
		.reset_in15     (1'b0),                                 // (terminated)
		.reset_req_in15 (1'b0)                                  // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (altpll_sys_c1_clk),                  //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_003 (
		.reset_in0      (~reset_reset_n),                       // reset_in0.reset
		.reset_in1      (nios2_gen2_debug_reset_request_reset), // reset_in1.reset
		.clk            (altpll_sys_c1_clk),                    //       clk.clk
		.reset_out      (rst_controller_003_reset_out_reset),   // reset_out.reset
		.reset_req      (),                                     // (terminated)
		.reset_req_in0  (1'b0),                                 // (terminated)
		.reset_req_in1  (1'b0),                                 // (terminated)
		.reset_in2      (1'b0),                                 // (terminated)
		.reset_req_in2  (1'b0),                                 // (terminated)
		.reset_in3      (1'b0),                                 // (terminated)
		.reset_req_in3  (1'b0),                                 // (terminated)
		.reset_in4      (1'b0),                                 // (terminated)
		.reset_req_in4  (1'b0),                                 // (terminated)
		.reset_in5      (1'b0),                                 // (terminated)
		.reset_req_in5  (1'b0),                                 // (terminated)
		.reset_in6      (1'b0),                                 // (terminated)
		.reset_req_in6  (1'b0),                                 // (terminated)
		.reset_in7      (1'b0),                                 // (terminated)
		.reset_req_in7  (1'b0),                                 // (terminated)
		.reset_in8      (1'b0),                                 // (terminated)
		.reset_req_in8  (1'b0),                                 // (terminated)
		.reset_in9      (1'b0),                                 // (terminated)
		.reset_req_in9  (1'b0),                                 // (terminated)
		.reset_in10     (1'b0),                                 // (terminated)
		.reset_req_in10 (1'b0),                                 // (terminated)
		.reset_in11     (1'b0),                                 // (terminated)
		.reset_req_in11 (1'b0),                                 // (terminated)
		.reset_in12     (1'b0),                                 // (terminated)
		.reset_req_in12 (1'b0),                                 // (terminated)
		.reset_in13     (1'b0),                                 // (terminated)
		.reset_req_in13 (1'b0),                                 // (terminated)
		.reset_in14     (1'b0),                                 // (terminated)
		.reset_req_in14 (1'b0),                                 // (terminated)
		.reset_in15     (1'b0),                                 // (terminated)
		.reset_req_in15 (1'b0)                                  // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_004 (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.clk            (clock_bridge_vip_out_clk_clk),           //       clk.clk
		.reset_out      (rst_controller_004_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_004_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_in1      (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_005 (
		.reset_in0      (nios2_gen2_debug_reset_request_reset), // reset_in0.reset
		.clk            (clk_clk),                              //       clk.clk
		.reset_out      (rst_controller_005_reset_out_reset),   // reset_out.reset
		.reset_req      (),                                     // (terminated)
		.reset_req_in0  (1'b0),                                 // (terminated)
		.reset_in1      (1'b0),                                 // (terminated)
		.reset_req_in1  (1'b0),                                 // (terminated)
		.reset_in2      (1'b0),                                 // (terminated)
		.reset_req_in2  (1'b0),                                 // (terminated)
		.reset_in3      (1'b0),                                 // (terminated)
		.reset_req_in3  (1'b0),                                 // (terminated)
		.reset_in4      (1'b0),                                 // (terminated)
		.reset_req_in4  (1'b0),                                 // (terminated)
		.reset_in5      (1'b0),                                 // (terminated)
		.reset_req_in5  (1'b0),                                 // (terminated)
		.reset_in6      (1'b0),                                 // (terminated)
		.reset_req_in6  (1'b0),                                 // (terminated)
		.reset_in7      (1'b0),                                 // (terminated)
		.reset_req_in7  (1'b0),                                 // (terminated)
		.reset_in8      (1'b0),                                 // (terminated)
		.reset_req_in8  (1'b0),                                 // (terminated)
		.reset_in9      (1'b0),                                 // (terminated)
		.reset_req_in9  (1'b0),                                 // (terminated)
		.reset_in10     (1'b0),                                 // (terminated)
		.reset_req_in10 (1'b0),                                 // (terminated)
		.reset_in11     (1'b0),                                 // (terminated)
		.reset_req_in11 (1'b0),                                 // (terminated)
		.reset_in12     (1'b0),                                 // (terminated)
		.reset_req_in12 (1'b0),                                 // (terminated)
		.reset_in13     (1'b0),                                 // (terminated)
		.reset_req_in13 (1'b0),                                 // (terminated)
		.reset_in14     (1'b0),                                 // (terminated)
		.reset_req_in14 (1'b0),                                 // (terminated)
		.reset_in15     (1'b0),                                 // (terminated)
		.reset_req_in15 (1'b0)                                  // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_006 (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.reset_in1      (nios2_gen2_debug_reset_request_reset),   // reset_in1.reset
		.clk            (clock_bridge_vip_out_clk_clk),           //       clk.clk
		.reset_out      (rst_controller_006_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_006_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_007 (
		.reset_in0      (nios2_gen2_debug_reset_request_reset), // reset_in0.reset
		.clk            (mem_if_ddr3_emif_afi_clk_clk),         //       clk.clk
		.reset_out      (rst_controller_007_reset_out_reset),   // reset_out.reset
		.reset_req      (),                                     // (terminated)
		.reset_req_in0  (1'b0),                                 // (terminated)
		.reset_in1      (1'b0),                                 // (terminated)
		.reset_req_in1  (1'b0),                                 // (terminated)
		.reset_in2      (1'b0),                                 // (terminated)
		.reset_req_in2  (1'b0),                                 // (terminated)
		.reset_in3      (1'b0),                                 // (terminated)
		.reset_req_in3  (1'b0),                                 // (terminated)
		.reset_in4      (1'b0),                                 // (terminated)
		.reset_req_in4  (1'b0),                                 // (terminated)
		.reset_in5      (1'b0),                                 // (terminated)
		.reset_req_in5  (1'b0),                                 // (terminated)
		.reset_in6      (1'b0),                                 // (terminated)
		.reset_req_in6  (1'b0),                                 // (terminated)
		.reset_in7      (1'b0),                                 // (terminated)
		.reset_req_in7  (1'b0),                                 // (terminated)
		.reset_in8      (1'b0),                                 // (terminated)
		.reset_req_in8  (1'b0),                                 // (terminated)
		.reset_in9      (1'b0),                                 // (terminated)
		.reset_req_in9  (1'b0),                                 // (terminated)
		.reset_in10     (1'b0),                                 // (terminated)
		.reset_req_in10 (1'b0),                                 // (terminated)
		.reset_in11     (1'b0),                                 // (terminated)
		.reset_req_in11 (1'b0),                                 // (terminated)
		.reset_in12     (1'b0),                                 // (terminated)
		.reset_req_in12 (1'b0),                                 // (terminated)
		.reset_in13     (1'b0),                                 // (terminated)
		.reset_req_in13 (1'b0),                                 // (terminated)
		.reset_in14     (1'b0),                                 // (terminated)
		.reset_req_in14 (1'b0),                                 // (terminated)
		.reset_in15     (1'b0),                                 // (terminated)
		.reset_req_in15 (1'b0)                                  // (terminated)
	);

endmodule
