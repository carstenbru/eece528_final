// megafunction wizard: %ALTSQRT%
// GENERATION: STANDARD
// VERSION: WM1.0
// MODULE: ALTSQRT 

// ============================================================
// File Name: sqrt.v
// Megafunction Name(s):
// 			ALTSQRT
//
// Simulation Library Files(s):
// 			altera_mf
// ============================================================
// ************************************************************
// THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
//
// 15.1.0 Build 185 10/21/2015 SJ Lite Edition
// ************************************************************


//Copyright (C) 1991-2015 Altera Corporation. All rights reserved.
//Your use of Altera Corporation's design tools, logic functions 
//and other software and tools, and its AMPP partner logic 
//functions, and any output files from any of the foregoing 
//(including device programming or simulation files), and any 
//associated documentation or information are expressly subject 
//to the terms and conditions of the Altera Program License 
//Subscription Agreement, the Altera Quartus Prime License Agreement,
//the Altera MegaCore Function License Agreement, or other 
//applicable license agreement, including, without limitation, 
//that your use is for the sole purpose of programming logic 
//devices manufactured by Altera and sold by Altera or its 
//authorized distributors.  Please refer to the applicable 
//agreement for further details.


// synopsys translate_off
`timescale 1 ps / 1 ps
// synopsys translate_on
module sqrt (
	clk,
	radical,
	q,
	remainder);

	input	  clk;
	input	[47:0]  radical;
	output	[23:0]  q;
	output	[24:0]  remainder;

	wire [23:0] sub_wire0;
	wire [24:0] sub_wire1;
	wire [23:0] q = sub_wire0[23:0];
	wire [24:0] remainder = sub_wire1[24:0];

	altsqrt	ALTSQRT_component (
				.clk (clk),
				.radical (radical),
				.q (sub_wire0),
				.remainder (sub_wire1)
				// synopsys translate_off
				,
				.aclr (),
				.ena ()
				// synopsys translate_on
				);
	defparam
		//ALTSQRT_component.pipeline = 2,
		ALTSQRT_component.q_port_width = 24,
		ALTSQRT_component.r_port_width = 25,
		ALTSQRT_component.width = 48;


endmodule

// ============================================================
// CNX file retrieval info
// ============================================================
// Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "MAX 10"
// Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
// Retrieval info: LIBRARY: altera_mf altera_mf.altera_mf_components.all
// Retrieval info: CONSTANT: PIPELINE NUMERIC "1"
// Retrieval info: CONSTANT: Q_PORT_WIDTH NUMERIC "24"
// Retrieval info: CONSTANT: R_PORT_WIDTH NUMERIC "25"
// Retrieval info: CONSTANT: WIDTH NUMERIC "48"
// Retrieval info: USED_PORT: clk 0 0 0 0 INPUT NODEFVAL "clk"
// Retrieval info: USED_PORT: q 0 0 24 0 OUTPUT NODEFVAL "q[23..0]"
// Retrieval info: USED_PORT: radical 0 0 48 0 INPUT NODEFVAL "radical[47..0]"
// Retrieval info: USED_PORT: remainder 0 0 25 0 OUTPUT NODEFVAL "remainder[24..0]"
// Retrieval info: CONNECT: @clk 0 0 0 0 clk 0 0 0 0
// Retrieval info: CONNECT: @radical 0 0 48 0 radical 0 0 48 0
// Retrieval info: CONNECT: q 0 0 24 0 @q 0 0 24 0
// Retrieval info: CONNECT: remainder 0 0 25 0 @remainder 0 0 25 0
// Retrieval info: GEN_FILE: TYPE_NORMAL sqrt.v TRUE
// Retrieval info: GEN_FILE: TYPE_NORMAL sqrt.inc FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL sqrt.cmp FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL sqrt.bsf FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL sqrt_inst.v FALSE
// Retrieval info: GEN_FILE: TYPE_NORMAL sqrt_bb.v FALSE
// Retrieval info: LIB_FILE: altera_mf
